reg [31:0] IMG_DATA [0:3071];

initial
begin
	IMG_DATA[0] = 32'h20201C;
	IMG_DATA[1] = 32'h403928;
	IMG_DATA[2] = 32'h342314;
	IMG_DATA[3] = 32'h342415;
	IMG_DATA[4] = 32'h352416;
	IMG_DATA[5] = 32'h362316;
	IMG_DATA[6] = 32'h3B2719;
	IMG_DATA[7] = 32'h382516;
	IMG_DATA[8] = 32'h3A2818;
	IMG_DATA[9] = 32'h3E2A1A;
	IMG_DATA[10] = 32'h3D2B19;
	IMG_DATA[11] = 32'h3E2A19;
	IMG_DATA[12] = 32'h3F2A1A;
	IMG_DATA[13] = 32'h3E2B1A;
	IMG_DATA[14] = 32'h3F2A19;
	IMG_DATA[15] = 32'h3F2A19;
	IMG_DATA[16] = 32'h3F2A19;
	IMG_DATA[17] = 32'h3F2B19;
	IMG_DATA[18] = 32'h402A19;
	IMG_DATA[19] = 32'h412A19;
	IMG_DATA[20] = 32'h432C1A;
	IMG_DATA[21] = 32'h442B1B;
	IMG_DATA[22] = 32'h432B1E;
	IMG_DATA[23] = 32'h422C1C;
	IMG_DATA[24] = 32'h422B1B;
	IMG_DATA[25] = 32'h432C1C;
	IMG_DATA[26] = 32'h432C1C;
	IMG_DATA[27] = 32'h432C1C;
	IMG_DATA[28] = 32'h432C1C;
	IMG_DATA[29] = 32'h432C1B;
	IMG_DATA[30] = 32'h422B1C;
	IMG_DATA[31] = 32'h422C1B;
	IMG_DATA[32] = 32'h432C1C;
	IMG_DATA[33] = 32'h432C1C;
	IMG_DATA[34] = 32'h422B1B;
	IMG_DATA[35] = 32'h432C1C;
	IMG_DATA[36] = 32'h432C1C;
	IMG_DATA[37] = 32'h442C1B;
	IMG_DATA[38] = 32'h432C1C;
	IMG_DATA[39] = 32'h432C1C;
	IMG_DATA[40] = 32'h442D1D;
	IMG_DATA[41] = 32'h432C1C;
	IMG_DATA[42] = 32'h432C1B;
	IMG_DATA[43] = 32'h432C1C;
	IMG_DATA[44] = 32'h432C1B;
	IMG_DATA[45] = 32'h432C1C;
	IMG_DATA[46] = 32'h432C1C;
	IMG_DATA[47] = 32'h432C1C;
	IMG_DATA[48] = 32'h432B1B;
	IMG_DATA[49] = 32'h442B1A;
	IMG_DATA[50] = 32'h422B1B;
	IMG_DATA[51] = 32'h442B1A;
	IMG_DATA[52] = 32'h412A1A;
	IMG_DATA[53] = 32'h422A1A;
	IMG_DATA[54] = 32'h412A19;
	IMG_DATA[55] = 32'h412A19;
	IMG_DATA[56] = 32'h402A1A;
	IMG_DATA[57] = 32'h3F2919;
	IMG_DATA[58] = 32'h402919;
	IMG_DATA[59] = 32'h402A19;
	IMG_DATA[60] = 32'h402A19;
	IMG_DATA[61] = 32'h3F2A18;
	IMG_DATA[62] = 32'h3F2B19;
	IMG_DATA[63] = 32'h3F2B19;
	IMG_DATA[64] = 32'h23211C;
	IMG_DATA[65] = 32'h413B28;
	IMG_DATA[66] = 32'h372415;
	IMG_DATA[67] = 32'h342214;
	IMG_DATA[68] = 32'h2F1E13;
	IMG_DATA[69] = 32'h382517;
	IMG_DATA[70] = 32'h382617;
	IMG_DATA[71] = 32'h352315;
	IMG_DATA[72] = 32'h3C2819;
	IMG_DATA[73] = 32'h3D291A;
	IMG_DATA[74] = 32'h3E2A19;
	IMG_DATA[75] = 32'h402A19;
	IMG_DATA[76] = 32'h3F2A1A;
	IMG_DATA[77] = 32'h402B1B;
	IMG_DATA[78] = 32'h402B19;
	IMG_DATA[79] = 32'h432A1A;
	IMG_DATA[80] = 32'h422B1A;
	IMG_DATA[81] = 32'h412B1A;
	IMG_DATA[82] = 32'h432B1B;
	IMG_DATA[83] = 32'h432B1B;
	IMG_DATA[84] = 32'h432B1B;
	IMG_DATA[85] = 32'h432B1B;
	IMG_DATA[86] = 32'h432C1D;
	IMG_DATA[87] = 32'h432C1C;
	IMG_DATA[88] = 32'h432C1C;
	IMG_DATA[89] = 32'h442D1D;
	IMG_DATA[90] = 32'h442D1D;
	IMG_DATA[91] = 32'h442D1D;
	IMG_DATA[92] = 32'h432E1D;
	IMG_DATA[93] = 32'h442E1E;
	IMG_DATA[94] = 32'h452E1E;
	IMG_DATA[95] = 32'h432E1E;
	IMG_DATA[96] = 32'h452F1E;
	IMG_DATA[97] = 32'h452E1E;
	IMG_DATA[98] = 32'h452E1E;
	IMG_DATA[99] = 32'h452F1E;
	IMG_DATA[100] = 32'h462F1F;
	IMG_DATA[101] = 32'h452E1E;
	IMG_DATA[102] = 32'h45301F;
	IMG_DATA[103] = 32'h452F1E;
	IMG_DATA[104] = 32'h442E1E;
	IMG_DATA[105] = 32'h452F1E;
	IMG_DATA[106] = 32'h442D1D;
	IMG_DATA[107] = 32'h442E1E;
	IMG_DATA[108] = 32'h442E1E;
	IMG_DATA[109] = 32'h432D1D;
	IMG_DATA[110] = 32'h432D1D;
	IMG_DATA[111] = 32'h432C1C;
	IMG_DATA[112] = 32'h412A1A;
	IMG_DATA[113] = 32'h432C1A;
	IMG_DATA[114] = 32'h432B1B;
	IMG_DATA[115] = 32'h432C1B;
	IMG_DATA[116] = 32'h422B1B;
	IMG_DATA[117] = 32'h432B1B;
	IMG_DATA[118] = 32'h422B1B;
	IMG_DATA[119] = 32'h422B1B;
	IMG_DATA[120] = 32'h432B1B;
	IMG_DATA[121] = 32'h402A19;
	IMG_DATA[122] = 32'h402A19;
	IMG_DATA[123] = 32'h422A19;
	IMG_DATA[124] = 32'h40291A;
	IMG_DATA[125] = 32'h412A19;
	IMG_DATA[126] = 32'h412A1A;
	IMG_DATA[127] = 32'h412A19;
	IMG_DATA[128] = 32'h2C2C22;
	IMG_DATA[129] = 32'h393527;
	IMG_DATA[130] = 32'h382719;
	IMG_DATA[131] = 32'h3D2618;
	IMG_DATA[132] = 32'h3B2518;
	IMG_DATA[133] = 32'h312116;
	IMG_DATA[134] = 32'h332013;
	IMG_DATA[135] = 32'h312013;
	IMG_DATA[136] = 32'h3A2516;
	IMG_DATA[137] = 32'h422B1A;
	IMG_DATA[138] = 32'h422B1B;
	IMG_DATA[139] = 32'h422C1C;
	IMG_DATA[140] = 32'h442D1D;
	IMG_DATA[141] = 32'h432C1C;
	IMG_DATA[142] = 32'h432D1C;
	IMG_DATA[143] = 32'h452D1D;
	IMG_DATA[144] = 32'h432C1C;
	IMG_DATA[145] = 32'h442E1E;
	IMG_DATA[146] = 32'h452E1E;
	IMG_DATA[147] = 32'h452E1E;
	IMG_DATA[148] = 32'h452E1E;
	IMG_DATA[149] = 32'h452E1F;
	IMG_DATA[150] = 32'h452E1E;
	IMG_DATA[151] = 32'h452E1E;
	IMG_DATA[152] = 32'h452E1E;
	IMG_DATA[153] = 32'h462F1F;
	IMG_DATA[154] = 32'h462E1E;
	IMG_DATA[155] = 32'h462F1F;
	IMG_DATA[156] = 32'h472F1E;
	IMG_DATA[157] = 32'h482F1F;
	IMG_DATA[158] = 32'h472F1F;
	IMG_DATA[159] = 32'h462F1F;
	IMG_DATA[160] = 32'h472F1F;
	IMG_DATA[161] = 32'h482E20;
	IMG_DATA[162] = 32'h482F20;
	IMG_DATA[163] = 32'h472F1F;
	IMG_DATA[164] = 32'h492F21;
	IMG_DATA[165] = 32'h482F1F;
	IMG_DATA[166] = 32'h48301F;
	IMG_DATA[167] = 32'h482F1F;
	IMG_DATA[168] = 32'h493020;
	IMG_DATA[169] = 32'h482F1F;
	IMG_DATA[170] = 32'h462F1F;
	IMG_DATA[171] = 32'h452E1F;
	IMG_DATA[172] = 32'h452F1F;
	IMG_DATA[173] = 32'h452E1E;
	IMG_DATA[174] = 32'h452F1F;
	IMG_DATA[175] = 32'h442E1E;
	IMG_DATA[176] = 32'h432E1D;
	IMG_DATA[177] = 32'h442D1D;
	IMG_DATA[178] = 32'h442D1D;
	IMG_DATA[179] = 32'h432D1D;
	IMG_DATA[180] = 32'h432C1C;
	IMG_DATA[181] = 32'h432C1C;
	IMG_DATA[182] = 32'h422C1B;
	IMG_DATA[183] = 32'h442C1C;
	IMG_DATA[184] = 32'h432C1B;
	IMG_DATA[185] = 32'h432C1B;
	IMG_DATA[186] = 32'h432B1C;
	IMG_DATA[187] = 32'h432C1B;
	IMG_DATA[188] = 32'h422C1C;
	IMG_DATA[189] = 32'h422B1B;
	IMG_DATA[190] = 32'h442B1B;
	IMG_DATA[191] = 32'h442C1A;
	IMG_DATA[192] = 32'h2B291F;
	IMG_DATA[193] = 32'h2A281D;
	IMG_DATA[194] = 32'h382A1D;
	IMG_DATA[195] = 32'h3F2A19;
	IMG_DATA[196] = 32'h422C1C;
	IMG_DATA[197] = 32'h362618;
	IMG_DATA[198] = 32'h261710;
	IMG_DATA[199] = 32'h2A1B12;
	IMG_DATA[200] = 32'h452D1D;
	IMG_DATA[201] = 32'h48301E;
	IMG_DATA[202] = 32'h49311E;
	IMG_DATA[203] = 32'h49321E;
	IMG_DATA[204] = 32'h49321D;
	IMG_DATA[205] = 32'h49321E;
	IMG_DATA[206] = 32'h4A331E;
	IMG_DATA[207] = 32'h493121;
	IMG_DATA[208] = 32'h493020;
	IMG_DATA[209] = 32'h493120;
	IMG_DATA[210] = 32'h48311E;
	IMG_DATA[211] = 32'h483120;
	IMG_DATA[212] = 32'h493120;
	IMG_DATA[213] = 32'h4A321F;
	IMG_DATA[214] = 32'h4A3120;
	IMG_DATA[215] = 32'h4A3121;
	IMG_DATA[216] = 32'h4A3120;
	IMG_DATA[217] = 32'h4B3221;
	IMG_DATA[218] = 32'h4A3120;
	IMG_DATA[219] = 32'h4B3221;
	IMG_DATA[220] = 32'h4C331F;
	IMG_DATA[221] = 32'h4A3120;
	IMG_DATA[222] = 32'h4B3220;
	IMG_DATA[223] = 32'h4A3321;
	IMG_DATA[224] = 32'h493121;
	IMG_DATA[225] = 32'h493020;
	IMG_DATA[226] = 32'h493020;
	IMG_DATA[227] = 32'h493121;
	IMG_DATA[228] = 32'h4A3122;
	IMG_DATA[229] = 32'h4A3121;
	IMG_DATA[230] = 32'h4A3121;
	IMG_DATA[231] = 32'h48311F;
	IMG_DATA[232] = 32'h4A3221;
	IMG_DATA[233] = 32'h4B3222;
	IMG_DATA[234] = 32'h4A3121;
	IMG_DATA[235] = 32'h483221;
	IMG_DATA[236] = 32'h473020;
	IMG_DATA[237] = 32'h483020;
	IMG_DATA[238] = 32'h48301E;
	IMG_DATA[239] = 32'h47301F;
	IMG_DATA[240] = 32'h472F1F;
	IMG_DATA[241] = 32'h472F1F;
	IMG_DATA[242] = 32'h472F1F;
	IMG_DATA[243] = 32'h483020;
	IMG_DATA[244] = 32'h472F1F;
	IMG_DATA[245] = 32'h472F1F;
	IMG_DATA[246] = 32'h452F1F;
	IMG_DATA[247] = 32'h462F1F;
	IMG_DATA[248] = 32'h452E1E;
	IMG_DATA[249] = 32'h452E1E;
	IMG_DATA[250] = 32'h452E1E;
	IMG_DATA[251] = 32'h442D1D;
	IMG_DATA[252] = 32'h442E1C;
	IMG_DATA[253] = 32'h422E1D;
	IMG_DATA[254] = 32'h422E1D;
	IMG_DATA[255] = 32'h442E1D;
	IMG_DATA[256] = 32'h27221A;
	IMG_DATA[257] = 32'h262118;
	IMG_DATA[258] = 32'h423826;
	IMG_DATA[259] = 32'h442D1C;
	IMG_DATA[260] = 32'h49311F;
	IMG_DATA[261] = 32'h493221;
	IMG_DATA[262] = 32'h2C2015;
	IMG_DATA[263] = 32'h271811;
	IMG_DATA[264] = 32'h513721;
	IMG_DATA[265] = 32'h503922;
	IMG_DATA[266] = 32'h4F3822;
	IMG_DATA[267] = 32'h503820;
	IMG_DATA[268] = 32'h503721;
	IMG_DATA[269] = 32'h4F3721;
	IMG_DATA[270] = 32'h4E3621;
	IMG_DATA[271] = 32'h4F3821;
	IMG_DATA[272] = 32'h503923;
	IMG_DATA[273] = 32'h513823;
	IMG_DATA[274] = 32'h513822;
	IMG_DATA[275] = 32'h4F3722;
	IMG_DATA[276] = 32'h503821;
	IMG_DATA[277] = 32'h503822;
	IMG_DATA[278] = 32'h503921;
	IMG_DATA[279] = 32'h4F3721;
	IMG_DATA[280] = 32'h4F3822;
	IMG_DATA[281] = 32'h513922;
	IMG_DATA[282] = 32'h513921;
	IMG_DATA[283] = 32'h4F3820;
	IMG_DATA[284] = 32'h503921;
	IMG_DATA[285] = 32'h503822;
	IMG_DATA[286] = 32'h4F3722;
	IMG_DATA[287] = 32'h4F3822;
	IMG_DATA[288] = 32'h4F3722;
	IMG_DATA[289] = 32'h4F3621;
	IMG_DATA[290] = 32'h4E3720;
	IMG_DATA[291] = 32'h4E3720;
	IMG_DATA[292] = 32'h4D3521;
	IMG_DATA[293] = 32'h4E3522;
	IMG_DATA[294] = 32'h4F3723;
	IMG_DATA[295] = 32'h4E3621;
	IMG_DATA[296] = 32'h4F3622;
	IMG_DATA[297] = 32'h4F3722;
	IMG_DATA[298] = 32'h4E3620;
	IMG_DATA[299] = 32'h4D3422;
	IMG_DATA[300] = 32'h4C3421;
	IMG_DATA[301] = 32'h4B3420;
	IMG_DATA[302] = 32'h4C3321;
	IMG_DATA[303] = 32'h4D3421;
	IMG_DATA[304] = 32'h4C3421;
	IMG_DATA[305] = 32'h4C3320;
	IMG_DATA[306] = 32'h4B3321;
	IMG_DATA[307] = 32'h4B3221;
	IMG_DATA[308] = 32'h493220;
	IMG_DATA[309] = 32'h493020;
	IMG_DATA[310] = 32'h483120;
	IMG_DATA[311] = 32'h49301E;
	IMG_DATA[312] = 32'h492F21;
	IMG_DATA[313] = 32'h49301F;
	IMG_DATA[314] = 32'h482F1F;
	IMG_DATA[315] = 32'h48301F;
	IMG_DATA[316] = 32'h452E1F;
	IMG_DATA[317] = 32'h462F1F;
	IMG_DATA[318] = 32'h462F1F;
	IMG_DATA[319] = 32'h462E1F;
	IMG_DATA[320] = 32'h2B2419;
	IMG_DATA[321] = 32'h2E2519;
	IMG_DATA[322] = 32'h433727;
	IMG_DATA[323] = 32'h453120;
	IMG_DATA[324] = 32'h4B331E;
	IMG_DATA[325] = 32'h503822;
	IMG_DATA[326] = 32'h42301F;
	IMG_DATA[327] = 32'h271A12;
	IMG_DATA[328] = 32'h583E27;
	IMG_DATA[329] = 32'h563C26;
	IMG_DATA[330] = 32'h563D25;
	IMG_DATA[331] = 32'h563D26;
	IMG_DATA[332] = 32'h583D25;
	IMG_DATA[333] = 32'h563C24;
	IMG_DATA[334] = 32'h563F26;
	IMG_DATA[335] = 32'h594027;
	IMG_DATA[336] = 32'h574026;
	IMG_DATA[337] = 32'h593E26;
	IMG_DATA[338] = 32'h583F26;
	IMG_DATA[339] = 32'h573E26;
	IMG_DATA[340] = 32'h553D26;
	IMG_DATA[341] = 32'h573C26;
	IMG_DATA[342] = 32'h563D25;
	IMG_DATA[343] = 32'h543C24;
	IMG_DATA[344] = 32'h573D25;
	IMG_DATA[345] = 32'h553D25;
	IMG_DATA[346] = 32'h563C25;
	IMG_DATA[347] = 32'h563D25;
	IMG_DATA[348] = 32'h563E25;
	IMG_DATA[349] = 32'h543D24;
	IMG_DATA[350] = 32'h553E26;
	IMG_DATA[351] = 32'h553D25;
	IMG_DATA[352] = 32'h553D25;
	IMG_DATA[353] = 32'h543D25;
	IMG_DATA[354] = 32'h533B24;
	IMG_DATA[355] = 32'h533C25;
	IMG_DATA[356] = 32'h553C26;
	IMG_DATA[357] = 32'h543B26;
	IMG_DATA[358] = 32'h543D26;
	IMG_DATA[359] = 32'h523A25;
	IMG_DATA[360] = 32'h523B25;
	IMG_DATA[361] = 32'h533B26;
	IMG_DATA[362] = 32'h513C2E;
	IMG_DATA[363] = 32'h503925;
	IMG_DATA[364] = 32'h5B4633;
	IMG_DATA[365] = 32'h513924;
	IMG_DATA[366] = 32'h503922;
	IMG_DATA[367] = 32'h503822;
	IMG_DATA[368] = 32'h4F3723;
	IMG_DATA[369] = 32'h4F3722;
	IMG_DATA[370] = 32'h4F3620;
	IMG_DATA[371] = 32'h4F3620;
	IMG_DATA[372] = 32'h4E3621;
	IMG_DATA[373] = 32'h4D3521;
	IMG_DATA[374] = 32'h4D3521;
	IMG_DATA[375] = 32'h4C3421;
	IMG_DATA[376] = 32'h4A331F;
	IMG_DATA[377] = 32'h4A331F;
	IMG_DATA[378] = 32'h4B3320;
	IMG_DATA[379] = 32'h4A3220;
	IMG_DATA[380] = 32'h4A3221;
	IMG_DATA[381] = 32'h493120;
	IMG_DATA[382] = 32'h493021;
	IMG_DATA[383] = 32'h4A3121;
	IMG_DATA[384] = 32'h34271A;
	IMG_DATA[385] = 32'h3F2B1D;
	IMG_DATA[386] = 32'h45301F;
	IMG_DATA[387] = 32'h4C3422;
	IMG_DATA[388] = 32'h58402F;
	IMG_DATA[389] = 32'h696564;
	IMG_DATA[390] = 32'h7D8FA1;
	IMG_DATA[391] = 32'h81A8C1;
	IMG_DATA[392] = 32'h86B1C5;
	IMG_DATA[393] = 32'h83A4B4;
	IMG_DATA[394] = 32'h767F81;
	IMG_DATA[395] = 32'h5C442F;
	IMG_DATA[396] = 32'h5E4329;
	IMG_DATA[397] = 32'h5E4229;
	IMG_DATA[398] = 32'h5E4329;
	IMG_DATA[399] = 32'h5E432A;
	IMG_DATA[400] = 32'h5C4328;
	IMG_DATA[401] = 32'h5E432A;
	IMG_DATA[402] = 32'h5D442A;
	IMG_DATA[403] = 32'h5F442B;
	IMG_DATA[404] = 32'h60462C;
	IMG_DATA[405] = 32'h5E442A;
	IMG_DATA[406] = 32'h5F442B;
	IMG_DATA[407] = 32'h5F442B;
	IMG_DATA[408] = 32'h5F432A;
	IMG_DATA[409] = 32'h5F432C;
	IMG_DATA[410] = 32'h5F442B;
	IMG_DATA[411] = 32'h60442B;
	IMG_DATA[412] = 32'h60452B;
	IMG_DATA[413] = 32'h5F452B;
	IMG_DATA[414] = 32'h5D452C;
	IMG_DATA[415] = 32'h5D442A;
	IMG_DATA[416] = 32'h5C4329;
	IMG_DATA[417] = 32'h5C432A;
	IMG_DATA[418] = 32'h5B4429;
	IMG_DATA[419] = 32'h5C422A;
	IMG_DATA[420] = 32'h5B432A;
	IMG_DATA[421] = 32'h5D4229;
	IMG_DATA[422] = 32'h594228;
	IMG_DATA[423] = 32'h5A4328;
	IMG_DATA[424] = 32'h604834;
	IMG_DATA[425] = 32'h604F47;
	IMG_DATA[426] = 32'h3B446D;
	IMG_DATA[427] = 32'h625E69;
	IMG_DATA[428] = 32'h999389;
	IMG_DATA[429] = 32'h604A37;
	IMG_DATA[430] = 32'h553D27;
	IMG_DATA[431] = 32'h543D27;
	IMG_DATA[432] = 32'h553D27;
	IMG_DATA[433] = 32'h543C27;
	IMG_DATA[434] = 32'h523B26;
	IMG_DATA[435] = 32'h523B24;
	IMG_DATA[436] = 32'h513A24;
	IMG_DATA[437] = 32'h513924;
	IMG_DATA[438] = 32'h503923;
	IMG_DATA[439] = 32'h503822;
	IMG_DATA[440] = 32'h4F3722;
	IMG_DATA[441] = 32'h503822;
	IMG_DATA[442] = 32'h503723;
	IMG_DATA[443] = 32'h4F3622;
	IMG_DATA[444] = 32'h4E3621;
	IMG_DATA[445] = 32'h4F3620;
	IMG_DATA[446] = 32'h4E3521;
	IMG_DATA[447] = 32'h4E3520;
	IMG_DATA[448] = 32'h593E27;
	IMG_DATA[449] = 32'h5B3F28;
	IMG_DATA[450] = 32'h5E432B;
	IMG_DATA[451] = 32'h72615C;
	IMG_DATA[452] = 32'h9BBDD6;
	IMG_DATA[453] = 32'hA4E2FD;
	IMG_DATA[454] = 32'h98E3FE;
	IMG_DATA[455] = 32'h8DE1FD;
	IMG_DATA[456] = 32'h83DDFC;
	IMG_DATA[457] = 32'h81DBFD;
	IMG_DATA[458] = 32'h80D9FC;
	IMG_DATA[459] = 32'h7DC6E4;
	IMG_DATA[460] = 32'h6D7167;
	IMG_DATA[461] = 32'h674C30;
	IMG_DATA[462] = 32'h654B2F;
	IMG_DATA[463] = 32'h654A2E;
	IMG_DATA[464] = 32'h654A2E;
	IMG_DATA[465] = 32'h654B2E;
	IMG_DATA[466] = 32'h65492E;
	IMG_DATA[467] = 32'h664B2F;
	IMG_DATA[468] = 32'h674C2F;
	IMG_DATA[469] = 32'h664C2F;
	IMG_DATA[470] = 32'h674D31;
	IMG_DATA[471] = 32'h664C2F;
	IMG_DATA[472] = 32'h664C30;
	IMG_DATA[473] = 32'h654B2E;
	IMG_DATA[474] = 32'h664C2E;
	IMG_DATA[475] = 32'h664C2E;
	IMG_DATA[476] = 32'h664C2F;
	IMG_DATA[477] = 32'h654A2E;
	IMG_DATA[478] = 32'h654A2E;
	IMG_DATA[479] = 32'h654A30;
	IMG_DATA[480] = 32'h654A2E;
	IMG_DATA[481] = 32'h63482E;
	IMG_DATA[482] = 32'h62482D;
	IMG_DATA[483] = 32'h61492D;
	IMG_DATA[484] = 32'h5F472C;
	IMG_DATA[485] = 32'h61452D;
	IMG_DATA[486] = 32'h62462D;
	IMG_DATA[487] = 32'h5F452D;
	IMG_DATA[488] = 32'h988F80;
	IMG_DATA[489] = 32'h847969;
	IMG_DATA[490] = 32'h4A5173;
	IMG_DATA[491] = 32'h494859;
	IMG_DATA[492] = 32'h644D39;
	IMG_DATA[493] = 32'h594329;
	IMG_DATA[494] = 32'h594228;
	IMG_DATA[495] = 32'h5A422A;
	IMG_DATA[496] = 32'h594229;
	IMG_DATA[497] = 32'h574127;
	IMG_DATA[498] = 32'h584128;
	IMG_DATA[499] = 32'h574026;
	IMG_DATA[500] = 32'h563F27;
	IMG_DATA[501] = 32'h573E27;
	IMG_DATA[502] = 32'h563D26;
	IMG_DATA[503] = 32'h563E26;
	IMG_DATA[504] = 32'h543D27;
	IMG_DATA[505] = 32'h533C26;
	IMG_DATA[506] = 32'h543D25;
	IMG_DATA[507] = 32'h523C25;
	IMG_DATA[508] = 32'h513A25;
	IMG_DATA[509] = 32'h523A25;
	IMG_DATA[510] = 32'h513A24;
	IMG_DATA[511] = 32'h513925;
	IMG_DATA[512] = 32'h66492D;
	IMG_DATA[513] = 32'h674B2E;
	IMG_DATA[514] = 32'h70605B;
	IMG_DATA[515] = 32'hA4CEEC;
	IMG_DATA[516] = 32'hAAE5FC;
	IMG_DATA[517] = 32'hA6E7FE;
	IMG_DATA[518] = 32'h98E3FD;
	IMG_DATA[519] = 32'h8FDFFE;
	IMG_DATA[520] = 32'h87DDFC;
	IMG_DATA[521] = 32'h83D9FD;
	IMG_DATA[522] = 32'h82DAFD;
	IMG_DATA[523] = 32'h7FDAFC;
	IMG_DATA[524] = 32'h7CD1F4;
	IMG_DATA[525] = 32'h727A72;
	IMG_DATA[526] = 32'h6C5031;
	IMG_DATA[527] = 32'h6D4F32;
	IMG_DATA[528] = 32'h6C4E30;
	IMG_DATA[529] = 32'h6D4F33;
	IMG_DATA[530] = 32'h6E5030;
	IMG_DATA[531] = 32'h6C4F31;
	IMG_DATA[532] = 32'h6B4E30;
	IMG_DATA[533] = 32'h6D5030;
	IMG_DATA[534] = 32'h6B4E30;
	IMG_DATA[535] = 32'h6B4E30;
	IMG_DATA[536] = 32'h6B4F2F;
	IMG_DATA[537] = 32'h6A4E30;
	IMG_DATA[538] = 32'h6A4D30;
	IMG_DATA[539] = 32'h6B4E30;
	IMG_DATA[540] = 32'h6B4E31;
	IMG_DATA[541] = 32'h694E31;
	IMG_DATA[542] = 32'h694D30;
	IMG_DATA[543] = 32'h684D31;
	IMG_DATA[544] = 32'h694E31;
	IMG_DATA[545] = 32'h694D32;
	IMG_DATA[546] = 32'h6B4E31;
	IMG_DATA[547] = 32'h694C31;
	IMG_DATA[548] = 32'h674C30;
	IMG_DATA[549] = 32'h674D30;
	IMG_DATA[550] = 32'h674A2F;
	IMG_DATA[551] = 32'h664B30;
	IMG_DATA[552] = 32'h674C30;
	IMG_DATA[553] = 32'h80715F;
	IMG_DATA[554] = 32'h64697F;
	IMG_DATA[555] = 32'h747B7D;
	IMG_DATA[556] = 32'h8C8478;
	IMG_DATA[557] = 32'h654D36;
	IMG_DATA[558] = 32'h60452D;
	IMG_DATA[559] = 32'h61432D;
	IMG_DATA[560] = 32'h5F432D;
	IMG_DATA[561] = 32'h5D442D;
	IMG_DATA[562] = 32'h5D442C;
	IMG_DATA[563] = 32'h5D432D;
	IMG_DATA[564] = 32'h5A442A;
	IMG_DATA[565] = 32'h5B442D;
	IMG_DATA[566] = 32'h5C412A;
	IMG_DATA[567] = 32'h5C432A;
	IMG_DATA[568] = 32'h5A4129;
	IMG_DATA[569] = 32'h5A4329;
	IMG_DATA[570] = 32'h5A4129;
	IMG_DATA[571] = 32'h5A4129;
	IMG_DATA[572] = 32'h594028;
	IMG_DATA[573] = 32'h5A3F29;
	IMG_DATA[574] = 32'h584028;
	IMG_DATA[575] = 32'h574029;
	IMG_DATA[576] = 32'h6F5232;
	IMG_DATA[577] = 32'h71563C;
	IMG_DATA[578] = 32'h95B8D6;
	IMG_DATA[579] = 32'hA5DFFD;
	IMG_DATA[580] = 32'hABE6FD;
	IMG_DATA[581] = 32'h9EE3FE;
	IMG_DATA[582] = 32'h8ADFFC;
	IMG_DATA[583] = 32'h83DBFC;
	IMG_DATA[584] = 32'h80D8FB;
	IMG_DATA[585] = 32'h87D9FD;
	IMG_DATA[586] = 32'h89DDFC;
	IMG_DATA[587] = 32'h81D7F8;
	IMG_DATA[588] = 32'h8FD3EC;
	IMG_DATA[589] = 32'hA7CBCF;
	IMG_DATA[590] = 32'hA0927A;
	IMG_DATA[591] = 32'h7D6344;
	IMG_DATA[592] = 32'h725435;
	IMG_DATA[593] = 32'h715535;
	IMG_DATA[594] = 32'h735534;
	IMG_DATA[595] = 32'h725534;
	IMG_DATA[596] = 32'h715533;
	IMG_DATA[597] = 32'h715434;
	IMG_DATA[598] = 32'h6F5333;
	IMG_DATA[599] = 32'h6E5232;
	IMG_DATA[600] = 32'h6F5332;
	IMG_DATA[601] = 32'h705433;
	IMG_DATA[602] = 32'h715535;
	IMG_DATA[603] = 32'h715434;
	IMG_DATA[604] = 32'h705332;
	IMG_DATA[605] = 32'h6F5333;
	IMG_DATA[606] = 32'h6E5132;
	IMG_DATA[607] = 32'h6F5132;
	IMG_DATA[608] = 32'h6F5232;
	IMG_DATA[609] = 32'h6D5131;
	IMG_DATA[610] = 32'h6D5031;
	IMG_DATA[611] = 32'h6D5032;
	IMG_DATA[612] = 32'h6D5032;
	IMG_DATA[613] = 32'h6F5134;
	IMG_DATA[614] = 32'h6F5233;
	IMG_DATA[615] = 32'h6D5032;
	IMG_DATA[616] = 32'h6B4F32;
	IMG_DATA[617] = 32'h76654E;
	IMG_DATA[618] = 32'h62534C;
	IMG_DATA[619] = 32'hBBC2BF;
	IMG_DATA[620] = 32'h70573F;
	IMG_DATA[621] = 32'h684C31;
	IMG_DATA[622] = 32'h654B30;
	IMG_DATA[623] = 32'h65492F;
	IMG_DATA[624] = 32'h664A30;
	IMG_DATA[625] = 32'h674A31;
	IMG_DATA[626] = 32'h664A31;
	IMG_DATA[627] = 32'h664A2F;
	IMG_DATA[628] = 32'h644831;
	IMG_DATA[629] = 32'h644730;
	IMG_DATA[630] = 32'h664930;
	IMG_DATA[631] = 32'h654830;
	IMG_DATA[632] = 32'h64482E;
	IMG_DATA[633] = 32'h63472E;
	IMG_DATA[634] = 32'h62452E;
	IMG_DATA[635] = 32'h61462F;
	IMG_DATA[636] = 32'h62452E;
	IMG_DATA[637] = 32'h60452E;
	IMG_DATA[638] = 32'h61462C;
	IMG_DATA[639] = 32'h60452D;
	IMG_DATA[640] = 32'h765836;
	IMG_DATA[641] = 32'h827672;
	IMG_DATA[642] = 32'h9DD8FC;
	IMG_DATA[643] = 32'hA2DEFD;
	IMG_DATA[644] = 32'hAFE4FD;
	IMG_DATA[645] = 32'hB0E3F4;
	IMG_DATA[646] = 32'hB4D4D8;
	IMG_DATA[647] = 32'hBACAC2;
	IMG_DATA[648] = 32'hB1C9C8;
	IMG_DATA[649] = 32'h9BD2E2;
	IMG_DATA[650] = 32'h79C7E8;
	IMG_DATA[651] = 32'hC4D7D8;
	IMG_DATA[652] = 32'hB4B5A1;
	IMG_DATA[653] = 32'h858576;
	IMG_DATA[654] = 32'h757669;
	IMG_DATA[655] = 32'hC5C4B3;
	IMG_DATA[656] = 32'h9A8668;
	IMG_DATA[657] = 32'h765937;
	IMG_DATA[658] = 32'h785837;
	IMG_DATA[659] = 32'h785837;
	IMG_DATA[660] = 32'h775937;
	IMG_DATA[661] = 32'h775837;
	IMG_DATA[662] = 32'h785938;
	IMG_DATA[663] = 32'h785938;
	IMG_DATA[664] = 32'h755837;
	IMG_DATA[665] = 32'h755938;
	IMG_DATA[666] = 32'h765837;
	IMG_DATA[667] = 32'h745736;
	IMG_DATA[668] = 32'h735635;
	IMG_DATA[669] = 32'h755635;
	IMG_DATA[670] = 32'h735535;
	IMG_DATA[671] = 32'h725535;
	IMG_DATA[672] = 32'h725535;
	IMG_DATA[673] = 32'h725534;
	IMG_DATA[674] = 32'h705435;
	IMG_DATA[675] = 32'h705434;
	IMG_DATA[676] = 32'h705434;
	IMG_DATA[677] = 32'h715433;
	IMG_DATA[678] = 32'h715535;
	IMG_DATA[679] = 32'h715434;
	IMG_DATA[680] = 32'h715437;
	IMG_DATA[681] = 32'h705436;
	IMG_DATA[682] = 32'h6F5434;
	IMG_DATA[683] = 32'hA5A298;
	IMG_DATA[684] = 32'h8F8170;
	IMG_DATA[685] = 32'h705235;
	IMG_DATA[686] = 32'h6F5135;
	IMG_DATA[687] = 32'h654B31;
	IMG_DATA[688] = 32'h56422D;
	IMG_DATA[689] = 32'h4B3A2C;
	IMG_DATA[690] = 32'h615247;
	IMG_DATA[691] = 32'h535453;
	IMG_DATA[692] = 32'h3F4144;
	IMG_DATA[693] = 32'h564738;
	IMG_DATA[694] = 32'h5B4532;
	IMG_DATA[695] = 32'h6A4F34;
	IMG_DATA[696] = 32'h684D32;
	IMG_DATA[697] = 32'h694D31;
	IMG_DATA[698] = 32'h674B31;
	IMG_DATA[699] = 32'h664C30;
	IMG_DATA[700] = 32'h674D2F;
	IMG_DATA[701] = 32'h684C31;
	IMG_DATA[702] = 32'h664C2E;
	IMG_DATA[703] = 32'h674D2F;
	IMG_DATA[704] = 32'h7C5D3A;
	IMG_DATA[705] = 32'h8A98A8;
	IMG_DATA[706] = 32'h93D7FB;
	IMG_DATA[707] = 32'hA3DEFC;
	IMG_DATA[708] = 32'hD2E9F3;
	IMG_DATA[709] = 32'hD9DBCC;
	IMG_DATA[710] = 32'h92927C;
	IMG_DATA[711] = 32'h5E6158;
	IMG_DATA[712] = 32'h686960;
	IMG_DATA[713] = 32'hA09E91;
	IMG_DATA[714] = 32'hCACDC3;
	IMG_DATA[715] = 32'hC2C3AC;
	IMG_DATA[716] = 32'h747261;
	IMG_DATA[717] = 32'h76776D;
	IMG_DATA[718] = 32'hADB1A1;
	IMG_DATA[719] = 32'h7D7F72;
	IMG_DATA[720] = 32'hC6C5B3;
	IMG_DATA[721] = 32'h876C49;
	IMG_DATA[722] = 32'h7A5C39;
	IMG_DATA[723] = 32'h7C5D3A;
	IMG_DATA[724] = 32'h7C5D3B;
	IMG_DATA[725] = 32'h7F5E3C;
	IMG_DATA[726] = 32'h7E5D3B;
	IMG_DATA[727] = 32'h7B5D3C;
	IMG_DATA[728] = 32'h795D3C;
	IMG_DATA[729] = 32'h7B5E3B;
	IMG_DATA[730] = 32'h795D3B;
	IMG_DATA[731] = 32'h785B3B;
	IMG_DATA[732] = 32'h785A3A;
	IMG_DATA[733] = 32'h795A3A;
	IMG_DATA[734] = 32'h7B5C3A;
	IMG_DATA[735] = 32'h7B5D3B;
	IMG_DATA[736] = 32'h7B5B3B;
	IMG_DATA[737] = 32'h775B3A;
	IMG_DATA[738] = 32'h785A3B;
	IMG_DATA[739] = 32'h765939;
	IMG_DATA[740] = 32'h745736;
	IMG_DATA[741] = 32'h745837;
	IMG_DATA[742] = 32'h745736;
	IMG_DATA[743] = 32'h755737;
	IMG_DATA[744] = 32'h745838;
	IMG_DATA[745] = 32'h725537;
	IMG_DATA[746] = 32'h725738;
	IMG_DATA[747] = 32'h968773;
	IMG_DATA[748] = 32'hBBBAB0;
	IMG_DATA[749] = 32'h6F5438;
	IMG_DATA[750] = 32'h584431;
	IMG_DATA[751] = 32'h474541;
	IMG_DATA[752] = 32'h5C788B;
	IMG_DATA[753] = 32'h7FB7D4;
	IMG_DATA[754] = 32'h91D4F6;
	IMG_DATA[755] = 32'h90D6F9;
	IMG_DATA[756] = 32'hABD2E0;
	IMG_DATA[757] = 32'hCBD2C6;
	IMG_DATA[758] = 32'hC6C4B4;
	IMG_DATA[759] = 32'hCFCEBE;
	IMG_DATA[760] = 32'hB0A794;
	IMG_DATA[761] = 32'h7B6148;
	IMG_DATA[762] = 32'h6B4F31;
	IMG_DATA[763] = 32'h6C4E32;
	IMG_DATA[764] = 32'h6A4F32;
	IMG_DATA[765] = 32'h6E5033;
	IMG_DATA[766] = 32'h6E5034;
	IMG_DATA[767] = 32'h6E5133;
	IMG_DATA[768] = 32'h846441;
	IMG_DATA[769] = 32'h8CABC0;
	IMG_DATA[770] = 32'h8BD4F7;
	IMG_DATA[771] = 32'hAFDFF3;
	IMG_DATA[772] = 32'hE8E8DD;
	IMG_DATA[773] = 32'h9FA18D;
	IMG_DATA[774] = 32'h858375;
	IMG_DATA[775] = 32'h888B81;
	IMG_DATA[776] = 32'h8D9190;
	IMG_DATA[777] = 32'hA2A898;
	IMG_DATA[778] = 32'hB7B7A4;
	IMG_DATA[779] = 32'h9EA08B;
	IMG_DATA[780] = 32'h999E89;
	IMG_DATA[781] = 32'h171B2A;
	IMG_DATA[782] = 32'h7B7B8B;
	IMG_DATA[783] = 32'hD0D8C5;
	IMG_DATA[784] = 32'hA1A197;
	IMG_DATA[785] = 32'hA79577;
	IMG_DATA[786] = 32'h81613E;
	IMG_DATA[787] = 32'h80603C;
	IMG_DATA[788] = 32'h80603C;
	IMG_DATA[789] = 32'h80603D;
	IMG_DATA[790] = 32'h80603B;
	IMG_DATA[791] = 32'h7F603D;
	IMG_DATA[792] = 32'h7D5F3D;
	IMG_DATA[793] = 32'h7B5E3C;
	IMG_DATA[794] = 32'h7E5E3C;
	IMG_DATA[795] = 32'h7E5E3C;
	IMG_DATA[796] = 32'h7E5E3B;
	IMG_DATA[797] = 32'h7F5F3B;
	IMG_DATA[798] = 32'h7F603C;
	IMG_DATA[799] = 32'h81603D;
	IMG_DATA[800] = 32'h7E5F3D;
	IMG_DATA[801] = 32'h7F603D;
	IMG_DATA[802] = 32'h80603C;
	IMG_DATA[803] = 32'h7E5F3C;
	IMG_DATA[804] = 32'h7B5C3B;
	IMG_DATA[805] = 32'h7A5C3B;
	IMG_DATA[806] = 32'h7A5D3B;
	IMG_DATA[807] = 32'h7A5D3B;
	IMG_DATA[808] = 32'h7A5D3C;
	IMG_DATA[809] = 32'h7A5B3A;
	IMG_DATA[810] = 32'h775A39;
	IMG_DATA[811] = 32'h765E3F;
	IMG_DATA[812] = 32'hC4CBC7;
	IMG_DATA[813] = 32'h675442;
	IMG_DATA[814] = 32'h6D7377;
	IMG_DATA[815] = 32'h97CEE9;
	IMG_DATA[816] = 32'h95DBF9;
	IMG_DATA[817] = 32'h98DBFA;
	IMG_DATA[818] = 32'h99DCF8;
	IMG_DATA[819] = 32'hC4DFDF;
	IMG_DATA[820] = 32'hBEC0B6;
	IMG_DATA[821] = 32'h4F525C;
	IMG_DATA[822] = 32'h2F3C4F;
	IMG_DATA[823] = 32'h4A5666;
	IMG_DATA[824] = 32'hB0B6AE;
	IMG_DATA[825] = 32'hD1CEBF;
	IMG_DATA[826] = 32'h7F674B;
	IMG_DATA[827] = 32'h715535;
	IMG_DATA[828] = 32'h715434;
	IMG_DATA[829] = 32'h6F5432;
	IMG_DATA[830] = 32'h725436;
	IMG_DATA[831] = 32'h705333;
	IMG_DATA[832] = 32'h866641;
	IMG_DATA[833] = 32'h88A7B9;
	IMG_DATA[834] = 32'h99CCDE;
	IMG_DATA[835] = 32'h99A195;
	IMG_DATA[836] = 32'hD7D7C2;
	IMG_DATA[837] = 32'h8A8B7E;
	IMG_DATA[838] = 32'hD4D6C4;
	IMG_DATA[839] = 32'h43494E;
	IMG_DATA[840] = 32'h333554;
	IMG_DATA[841] = 32'hD7DBCD;
	IMG_DATA[842] = 32'hA3A698;
	IMG_DATA[843] = 32'h9EA08E;
	IMG_DATA[844] = 32'hDADCCB;
	IMG_DATA[845] = 32'h888D92;
	IMG_DATA[846] = 32'hB3B3B2;
	IMG_DATA[847] = 32'hD6DECC;
	IMG_DATA[848] = 32'hA6A79A;
	IMG_DATA[849] = 32'hA8997C;
	IMG_DATA[850] = 32'h866542;
	IMG_DATA[851] = 32'h846340;
	IMG_DATA[852] = 32'h836340;
	IMG_DATA[853] = 32'h846240;
	IMG_DATA[854] = 32'h836340;
	IMG_DATA[855] = 32'h82623F;
	IMG_DATA[856] = 32'h82623F;
	IMG_DATA[857] = 32'h836542;
	IMG_DATA[858] = 32'h8B6D4F;
	IMG_DATA[859] = 32'h93816E;
	IMG_DATA[860] = 32'h988E81;
	IMG_DATA[861] = 32'h948879;
	IMG_DATA[862] = 32'h8E785F;
	IMG_DATA[863] = 32'hA08E75;
	IMG_DATA[864] = 32'hB9B199;
	IMG_DATA[865] = 32'hB4A991;
	IMG_DATA[866] = 32'h927659;
	IMG_DATA[867] = 32'h7F603E;
	IMG_DATA[868] = 32'h7C5F3C;
	IMG_DATA[869] = 32'h7F5F3C;
	IMG_DATA[870] = 32'h7F603D;
	IMG_DATA[871] = 32'h80603D;
	IMG_DATA[872] = 32'h7D5F3D;
	IMG_DATA[873] = 32'h7C5E3D;
	IMG_DATA[874] = 32'h785B3C;
	IMG_DATA[875] = 32'h7A5B3C;
	IMG_DATA[876] = 32'hA09F96;
	IMG_DATA[877] = 32'h98B4BF;
	IMG_DATA[878] = 32'h9CDAF3;
	IMG_DATA[879] = 32'h9CDEFB;
	IMG_DATA[880] = 32'h9CDEFB;
	IMG_DATA[881] = 32'hAAE1FA;
	IMG_DATA[882] = 32'hB4D7E5;
	IMG_DATA[883] = 32'hECEDE8;
	IMG_DATA[884] = 32'h6F7477;
	IMG_DATA[885] = 32'h8C9692;
	IMG_DATA[886] = 32'h818C8B;
	IMG_DATA[887] = 32'hABB8B6;
	IMG_DATA[888] = 32'h6F7E90;
	IMG_DATA[889] = 32'hC2C6BD;
	IMG_DATA[890] = 32'hC6BBAD;
	IMG_DATA[891] = 32'h785B3B;
	IMG_DATA[892] = 32'h765839;
	IMG_DATA[893] = 32'h765736;
	IMG_DATA[894] = 32'h765838;
	IMG_DATA[895] = 32'h745737;
	IMG_DATA[896] = 32'h896A44;
	IMG_DATA[897] = 32'h888065;
	IMG_DATA[898] = 32'h787561;
	IMG_DATA[899] = 32'h948F7B;
	IMG_DATA[900] = 32'hC9C8B1;
	IMG_DATA[901] = 32'h9B9C8F;
	IMG_DATA[902] = 32'hE2E4D5;
	IMG_DATA[903] = 32'hCCD0C1;
	IMG_DATA[904] = 32'hC0C2BF;
	IMG_DATA[905] = 32'hD6DECC;
	IMG_DATA[906] = 32'hB1B5A6;
	IMG_DATA[907] = 32'hBEC0AD;
	IMG_DATA[908] = 32'hCBCEC0;
	IMG_DATA[909] = 32'hE8ECD9;
	IMG_DATA[910] = 32'hE2E8D5;
	IMG_DATA[911] = 32'hC0C8B9;
	IMG_DATA[912] = 32'hC1BEAE;
	IMG_DATA[913] = 32'h9C8664;
	IMG_DATA[914] = 32'h886844;
	IMG_DATA[915] = 32'h886843;
	IMG_DATA[916] = 32'h896A43;
	IMG_DATA[917] = 32'h8A6B43;
	IMG_DATA[918] = 32'h8A6B45;
	IMG_DATA[919] = 32'h896A47;
	IMG_DATA[920] = 32'hA08C72;
	IMG_DATA[921] = 32'hCBC3AE;
	IMG_DATA[922] = 32'hC0BFAF;
	IMG_DATA[923] = 32'hC6CABB;
	IMG_DATA[924] = 32'hC8DAD6;
	IMG_DATA[925] = 32'hB5E1F5;
	IMG_DATA[926] = 32'hDFEAE3;
	IMG_DATA[927] = 32'hA3A69C;
	IMG_DATA[928] = 32'h727675;
	IMG_DATA[929] = 32'h7F8683;
	IMG_DATA[930] = 32'hC9C9BA;
	IMG_DATA[931] = 32'h9F8B6E;
	IMG_DATA[932] = 32'h816240;
	IMG_DATA[933] = 32'h81613E;
	IMG_DATA[934] = 32'h82623F;
	IMG_DATA[935] = 32'h81613E;
	IMG_DATA[936] = 32'h80603E;
	IMG_DATA[937] = 32'h80603E;
	IMG_DATA[938] = 32'h82613F;
	IMG_DATA[939] = 32'h7F613F;
	IMG_DATA[940] = 32'h868B87;
	IMG_DATA[941] = 32'hA1DBF6;
	IMG_DATA[942] = 32'h9DDFFA;
	IMG_DATA[943] = 32'h9CDFFA;
	IMG_DATA[944] = 32'hA4DFFB;
	IMG_DATA[945] = 32'hB0DCF4;
	IMG_DATA[946] = 32'hDFE6E2;
	IMG_DATA[947] = 32'hD8D9D2;
	IMG_DATA[948] = 32'hA1AA9B;
	IMG_DATA[949] = 32'h747A83;
	IMG_DATA[950] = 32'h181F37;
	IMG_DATA[951] = 32'h515C76;
	IMG_DATA[952] = 32'hD9E1D2;
	IMG_DATA[953] = 32'h8F9493;
	IMG_DATA[954] = 32'hDEDED1;
	IMG_DATA[955] = 32'h8A6F53;
	IMG_DATA[956] = 32'h7C5E3C;
	IMG_DATA[957] = 32'h785B3C;
	IMG_DATA[958] = 32'h775A3B;
	IMG_DATA[959] = 32'h775B3B;
	IMG_DATA[960] = 32'h8D6D44;
	IMG_DATA[961] = 32'h887B5A;
	IMG_DATA[962] = 32'h636D5F;
	IMG_DATA[963] = 32'h86846F;
	IMG_DATA[964] = 32'hABA48D;
	IMG_DATA[965] = 32'hB5B6A1;
	IMG_DATA[966] = 32'hCCD0C5;
	IMG_DATA[967] = 32'hE3E9D8;
	IMG_DATA[968] = 32'hDCE4D3;
	IMG_DATA[969] = 32'hBDC6BB;
	IMG_DATA[970] = 32'hC8C7B6;
	IMG_DATA[971] = 32'hB6B39A;
	IMG_DATA[972] = 32'hC4C7B5;
	IMG_DATA[973] = 32'hB9CBCB;
	IMG_DATA[974] = 32'hA3BCC1;
	IMG_DATA[975] = 32'h9EAAAA;
	IMG_DATA[976] = 32'hBAAF91;
	IMG_DATA[977] = 32'h92734C;
	IMG_DATA[978] = 32'h8E7047;
	IMG_DATA[979] = 32'h8E6F46;
	IMG_DATA[980] = 32'h8D6F46;
	IMG_DATA[981] = 32'h8D6E46;
	IMG_DATA[982] = 32'h907251;
	IMG_DATA[983] = 32'hB3B4B5;
	IMG_DATA[984] = 32'hE9EAE3;
	IMG_DATA[985] = 32'h7F857D;
	IMG_DATA[986] = 32'h828987;
	IMG_DATA[987] = 32'h929A96;
	IMG_DATA[988] = 32'hA1A59B;
	IMG_DATA[989] = 32'hD6DAC9;
	IMG_DATA[990] = 32'hB6B8A8;
	IMG_DATA[991] = 32'hAFB3A7;
	IMG_DATA[992] = 32'hC2CAB9;
	IMG_DATA[993] = 32'hECF2E0;
	IMG_DATA[994] = 32'hAAAFA5;
	IMG_DATA[995] = 32'hD0CFBE;
	IMG_DATA[996] = 32'h8B6A49;
	IMG_DATA[997] = 32'h896845;
	IMG_DATA[998] = 32'h866542;
	IMG_DATA[999] = 32'h84623F;
	IMG_DATA[1000] = 32'h856542;
	IMG_DATA[1001] = 32'h856441;
	IMG_DATA[1002] = 32'h866644;
	IMG_DATA[1003] = 32'h846A4B;
	IMG_DATA[1004] = 32'h98C3D5;
	IMG_DATA[1005] = 32'h96DAF8;
	IMG_DATA[1006] = 32'h96DCF9;
	IMG_DATA[1007] = 32'h95DDF9;
	IMG_DATA[1008] = 32'hA8E1F9;
	IMG_DATA[1009] = 32'hA7C8D8;
	IMG_DATA[1010] = 32'hD2D8D3;
	IMG_DATA[1011] = 32'hD7D9D0;
	IMG_DATA[1012] = 32'hCFD6C5;
	IMG_DATA[1013] = 32'h9DA1A6;
	IMG_DATA[1014] = 32'h212741;
	IMG_DATA[1015] = 32'h47506E;
	IMG_DATA[1016] = 32'hE2E9D8;
	IMG_DATA[1017] = 32'hA8ACA5;
	IMG_DATA[1018] = 32'hD4D7C9;
	IMG_DATA[1019] = 32'hA18B74;
	IMG_DATA[1020] = 32'h7E603D;
	IMG_DATA[1021] = 32'h7E5F3C;
	IMG_DATA[1022] = 32'h7C5F3D;
	IMG_DATA[1023] = 32'h7C5F3C;
	IMG_DATA[1024] = 32'h917249;
	IMG_DATA[1025] = 32'h91816D;
	IMG_DATA[1026] = 32'h7AC5E2;
	IMG_DATA[1027] = 32'h65A9C0;
	IMG_DATA[1028] = 32'h7C918D;
	IMG_DATA[1029] = 32'hB1AD9B;
	IMG_DATA[1030] = 32'hBEC2B1;
	IMG_DATA[1031] = 32'hB2C6C8;
	IMG_DATA[1032] = 32'h9FBCC4;
	IMG_DATA[1033] = 32'hADB4B0;
	IMG_DATA[1034] = 32'h9D9C8C;
	IMG_DATA[1035] = 32'h212734;
	IMG_DATA[1036] = 32'h79776C;
	IMG_DATA[1037] = 32'hB4B19C;
	IMG_DATA[1038] = 32'hB2B2A3;
	IMG_DATA[1039] = 32'h9C9E8D;
	IMG_DATA[1040] = 32'h957753;
	IMG_DATA[1041] = 32'h93704A;
	IMG_DATA[1042] = 32'h93714B;
	IMG_DATA[1043] = 32'h93714B;
	IMG_DATA[1044] = 32'h8F7048;
	IMG_DATA[1045] = 32'h8E6E4B;
	IMG_DATA[1046] = 32'hA5AEAC;
	IMG_DATA[1047] = 32'hD5EBF1;
	IMG_DATA[1048] = 32'hBEBFB2;
	IMG_DATA[1049] = 32'hC0C5B7;
	IMG_DATA[1050] = 32'hCCD0C4;
	IMG_DATA[1051] = 32'h6E7785;
	IMG_DATA[1052] = 32'hDAE0D1;
	IMG_DATA[1053] = 32'hC9C9BC;
	IMG_DATA[1054] = 32'hB2B6A4;
	IMG_DATA[1055] = 32'hD3DAC9;
	IMG_DATA[1056] = 32'h223C39;
	IMG_DATA[1057] = 32'h98AFA1;
	IMG_DATA[1058] = 32'hE6ECDC;
	IMG_DATA[1059] = 32'hC0C2B4;
	IMG_DATA[1060] = 32'h9E8667;
	IMG_DATA[1061] = 32'h8A6A44;
	IMG_DATA[1062] = 32'h8A6846;
	IMG_DATA[1063] = 32'h886744;
	IMG_DATA[1064] = 32'h896645;
	IMG_DATA[1065] = 32'h8A6845;
	IMG_DATA[1066] = 32'h8A6946;
	IMG_DATA[1067] = 32'h847B6A;
	IMG_DATA[1068] = 32'h83D0F2;
	IMG_DATA[1069] = 32'h82D7F6;
	IMG_DATA[1070] = 32'h86D6F5;
	IMG_DATA[1071] = 32'h74B2CB;
	IMG_DATA[1072] = 32'h6B868D;
	IMG_DATA[1073] = 32'h898C7F;
	IMG_DATA[1074] = 32'h9EA193;
	IMG_DATA[1075] = 32'hEAEADF;
	IMG_DATA[1076] = 32'hD7DCCC;
	IMG_DATA[1077] = 32'hEFF3E2;
	IMG_DATA[1078] = 32'hBFC2BA;
	IMG_DATA[1079] = 32'hCCD2C3;
	IMG_DATA[1080] = 32'hE4E8D9;
	IMG_DATA[1081] = 32'hB8BFB5;
	IMG_DATA[1082] = 32'hD4D5CA;
	IMG_DATA[1083] = 32'h9D886F;
	IMG_DATA[1084] = 32'h836442;
	IMG_DATA[1085] = 32'h836442;
	IMG_DATA[1086] = 32'h836340;
	IMG_DATA[1087] = 32'h846340;
	IMG_DATA[1088] = 32'h95764C;
	IMG_DATA[1089] = 32'h947B5E;
	IMG_DATA[1090] = 32'h8ACFED;
	IMG_DATA[1091] = 32'h74CCED;
	IMG_DATA[1092] = 32'h6AC4E5;
	IMG_DATA[1093] = 32'h6298AE;
	IMG_DATA[1094] = 32'h7B837F;
	IMG_DATA[1095] = 32'h9C998A;
	IMG_DATA[1096] = 32'hA4A597;
	IMG_DATA[1097] = 32'h757E7B;
	IMG_DATA[1098] = 32'h20415F;
	IMG_DATA[1099] = 32'h133D65;
	IMG_DATA[1100] = 32'h1C4B73;
	IMG_DATA[1101] = 32'h224A6A;
	IMG_DATA[1102] = 32'h2D5777;
	IMG_DATA[1103] = 32'h376687;
	IMG_DATA[1104] = 32'h896E4E;
	IMG_DATA[1105] = 32'h91714A;
	IMG_DATA[1106] = 32'h92704A;
	IMG_DATA[1107] = 32'h91714B;
	IMG_DATA[1108] = 32'h927149;
	IMG_DATA[1109] = 32'h958875;
	IMG_DATA[1110] = 32'hBFD2CE;
	IMG_DATA[1111] = 32'hC2C6BF;
	IMG_DATA[1112] = 32'hBDC0B1;
	IMG_DATA[1113] = 32'hEFF3E3;
	IMG_DATA[1114] = 32'hB8BFB7;
	IMG_DATA[1115] = 32'h313B58;
	IMG_DATA[1116] = 32'hC2C8C2;
	IMG_DATA[1117] = 32'hCCD0C3;
	IMG_DATA[1118] = 32'hCACDBD;
	IMG_DATA[1119] = 32'hF4F9E8;
	IMG_DATA[1120] = 32'hA6B6A7;
	IMG_DATA[1121] = 32'hDEE8D5;
	IMG_DATA[1122] = 32'hE7EFDD;
	IMG_DATA[1123] = 32'hCFD1C3;
	IMG_DATA[1124] = 32'h9D8568;
	IMG_DATA[1125] = 32'h8B6846;
	IMG_DATA[1126] = 32'h8A6745;
	IMG_DATA[1127] = 32'h896745;
	IMG_DATA[1128] = 32'h886745;
	IMG_DATA[1129] = 32'h8B6946;
	IMG_DATA[1130] = 32'h8C6B46;
	IMG_DATA[1131] = 32'h778986;
	IMG_DATA[1132] = 32'h66C2E2;
	IMG_DATA[1133] = 32'h5F9DB5;
	IMG_DATA[1134] = 32'h32474F;
	IMG_DATA[1135] = 32'h292E2C;
	IMG_DATA[1136] = 32'h323531;
	IMG_DATA[1137] = 32'h828277;
	IMG_DATA[1138] = 32'h686F6B;
	IMG_DATA[1139] = 32'hCBCCBD;
	IMG_DATA[1140] = 32'hDADECE;
	IMG_DATA[1141] = 32'hE8ECDB;
	IMG_DATA[1142] = 32'hE7EEDB;
	IMG_DATA[1143] = 32'hE5EBD9;
	IMG_DATA[1144] = 32'hD8DFD1;
	IMG_DATA[1145] = 32'hBAC1BB;
	IMG_DATA[1146] = 32'hD1D2C5;
	IMG_DATA[1147] = 32'h7B6654;
	IMG_DATA[1148] = 32'h846340;
	IMG_DATA[1149] = 32'h876744;
	IMG_DATA[1150] = 32'h8A6846;
	IMG_DATA[1151] = 32'h876743;
	IMG_DATA[1152] = 32'h95754D;
	IMG_DATA[1153] = 32'h967552;
	IMG_DATA[1154] = 32'h8BC3E0;
	IMG_DATA[1155] = 32'h7CD3F3;
	IMG_DATA[1156] = 32'h7CD3F4;
	IMG_DATA[1157] = 32'h70CAEB;
	IMG_DATA[1158] = 32'h53AACC;
	IMG_DATA[1159] = 32'h32779C;
	IMG_DATA[1160] = 32'h1F577D;
	IMG_DATA[1161] = 32'h1B547C;
	IMG_DATA[1162] = 32'h22628A;
	IMG_DATA[1163] = 32'h307EA9;
	IMG_DATA[1164] = 32'h3C95BF;
	IMG_DATA[1165] = 32'h3A8EB5;
	IMG_DATA[1166] = 32'h367DA4;
	IMG_DATA[1167] = 32'h356F93;
	IMG_DATA[1168] = 32'h806D55;
	IMG_DATA[1169] = 32'h93724B;
	IMG_DATA[1170] = 32'h96744E;
	IMG_DATA[1171] = 32'h93744D;
	IMG_DATA[1172] = 32'h95754D;
	IMG_DATA[1173] = 32'h8E938A;
	IMG_DATA[1174] = 32'h7F8072;
	IMG_DATA[1175] = 32'h888578;
	IMG_DATA[1176] = 32'hDCDDCE;
	IMG_DATA[1177] = 32'hE9EFDE;
	IMG_DATA[1178] = 32'hF9FCE9;
	IMG_DATA[1179] = 32'hECEEDE;
	IMG_DATA[1180] = 32'hEFF3E1;
	IMG_DATA[1181] = 32'hDBDCCE;
	IMG_DATA[1182] = 32'hD2D3C0;
	IMG_DATA[1183] = 32'hE5E9D8;
	IMG_DATA[1184] = 32'hF2F6E4;
	IMG_DATA[1185] = 32'hECF2E0;
	IMG_DATA[1186] = 32'hD9DDCD;
	IMG_DATA[1187] = 32'hC7C3AF;
	IMG_DATA[1188] = 32'h8E704E;
	IMG_DATA[1189] = 32'h8C6948;
	IMG_DATA[1190] = 32'h8D6A48;
	IMG_DATA[1191] = 32'h8C6A47;
	IMG_DATA[1192] = 32'h8C6948;
	IMG_DATA[1193] = 32'h8C6B48;
	IMG_DATA[1194] = 32'h8F6D47;
	IMG_DATA[1195] = 32'h656963;
	IMG_DATA[1196] = 32'h253841;
	IMG_DATA[1197] = 32'h1C2022;
	IMG_DATA[1198] = 32'h22292C;
	IMG_DATA[1199] = 32'h253B48;
	IMG_DATA[1200] = 32'h315970;
	IMG_DATA[1201] = 32'h678495;
	IMG_DATA[1202] = 32'h708899;
	IMG_DATA[1203] = 32'h989F9D;
	IMG_DATA[1204] = 32'hD2D2C0;
	IMG_DATA[1205] = 32'hD7DBCB;
	IMG_DATA[1206] = 32'hD7DFD1;
	IMG_DATA[1207] = 32'hCDD9D0;
	IMG_DATA[1208] = 32'hA9BDC2;
	IMG_DATA[1209] = 32'hB7BCB7;
	IMG_DATA[1210] = 32'h9BA49F;
	IMG_DATA[1211] = 32'h656D72;
	IMG_DATA[1212] = 32'h8A6945;
	IMG_DATA[1213] = 32'h896745;
	IMG_DATA[1214] = 32'h896845;
	IMG_DATA[1215] = 32'h8B6846;
	IMG_DATA[1216] = 32'h94754E;
	IMG_DATA[1217] = 32'h997751;
	IMG_DATA[1218] = 32'h8DB9CF;
	IMG_DATA[1219] = 32'h80D4F5;
	IMG_DATA[1220] = 32'h82D6F7;
	IMG_DATA[1221] = 32'h80D5F5;
	IMG_DATA[1222] = 32'h79CFEF;
	IMG_DATA[1223] = 32'h6AC1DF;
	IMG_DATA[1224] = 32'h59B0D0;
	IMG_DATA[1225] = 32'h4BA2C5;
	IMG_DATA[1226] = 32'h4AA8CD;
	IMG_DATA[1227] = 32'h50B1D8;
	IMG_DATA[1228] = 32'h54B4DC;
	IMG_DATA[1229] = 32'h51B2D7;
	IMG_DATA[1230] = 32'h459EC3;
	IMG_DATA[1231] = 32'h3B83A9;
	IMG_DATA[1232] = 32'h776F61;
	IMG_DATA[1233] = 32'h96744D;
	IMG_DATA[1234] = 32'h93714A;
	IMG_DATA[1235] = 32'h95744D;
	IMG_DATA[1236] = 32'h93724D;
	IMG_DATA[1237] = 32'h5C533C;
	IMG_DATA[1238] = 32'h56554D;
	IMG_DATA[1239] = 32'h767463;
	IMG_DATA[1240] = 32'hBCB9A8;
	IMG_DATA[1241] = 32'hD8DCCB;
	IMG_DATA[1242] = 32'hE9EDDD;
	IMG_DATA[1243] = 32'hE8EEDD;
	IMG_DATA[1244] = 32'hDCE3D2;
	IMG_DATA[1245] = 32'hC5C7B6;
	IMG_DATA[1246] = 32'h65665B;
	IMG_DATA[1247] = 32'hC3C5B3;
	IMG_DATA[1248] = 32'hD6D9C7;
	IMG_DATA[1249] = 32'hD4D4C4;
	IMG_DATA[1250] = 32'hB9BAA5;
	IMG_DATA[1251] = 32'h867D6D;
	IMG_DATA[1252] = 32'h8F6E4B;
	IMG_DATA[1253] = 32'h8C6C48;
	IMG_DATA[1254] = 32'h8B6B48;
	IMG_DATA[1255] = 32'h8B6A48;
	IMG_DATA[1256] = 32'h8F6D49;
	IMG_DATA[1257] = 32'h8F6D49;
	IMG_DATA[1258] = 32'h916E48;
	IMG_DATA[1259] = 32'h564432;
	IMG_DATA[1260] = 32'h162630;
	IMG_DATA[1261] = 32'h2A5E79;
	IMG_DATA[1262] = 32'h4EA2C7;
	IMG_DATA[1263] = 32'h67C3E8;
	IMG_DATA[1264] = 32'h7ED3F4;
	IMG_DATA[1265] = 32'h97D7F2;
	IMG_DATA[1266] = 32'h86BCDB;
	IMG_DATA[1267] = 32'h8EACC3;
	IMG_DATA[1268] = 32'h98A09E;
	IMG_DATA[1269] = 32'hBCBAA8;
	IMG_DATA[1270] = 32'hC7C8B2;
	IMG_DATA[1271] = 32'hC5C7B9;
	IMG_DATA[1272] = 32'hC0BFAE;
	IMG_DATA[1273] = 32'h9BA194;
	IMG_DATA[1274] = 32'h396C8B;
	IMG_DATA[1275] = 32'h4E7289;
	IMG_DATA[1276] = 32'h8A6745;
	IMG_DATA[1277] = 32'h876745;
	IMG_DATA[1278] = 32'h896845;
	IMG_DATA[1279] = 32'h886845;
	IMG_DATA[1280] = 32'h997851;
	IMG_DATA[1281] = 32'h997952;
	IMG_DATA[1282] = 32'h90AAB7;
	IMG_DATA[1283] = 32'h80D3F5;
	IMG_DATA[1284] = 32'h86D8F8;
	IMG_DATA[1285] = 32'h85D8F8;
	IMG_DATA[1286] = 32'h89D7F7;
	IMG_DATA[1287] = 32'h8CD5F5;
	IMG_DATA[1288] = 32'h89D4F0;
	IMG_DATA[1289] = 32'h7CCFEC;
	IMG_DATA[1290] = 32'h6DC7EB;
	IMG_DATA[1291] = 32'h65C5E9;
	IMG_DATA[1292] = 32'h61C2E7;
	IMG_DATA[1293] = 32'h5CBBE1;
	IMG_DATA[1294] = 32'h4FADD1;
	IMG_DATA[1295] = 32'h4091B5;
	IMG_DATA[1296] = 32'h6D726D;
	IMG_DATA[1297] = 32'h9C7C51;
	IMG_DATA[1298] = 32'h9B7B53;
	IMG_DATA[1299] = 32'h987651;
	IMG_DATA[1300] = 32'h8D704D;
	IMG_DATA[1301] = 32'h436975;
	IMG_DATA[1302] = 32'h468CAC;
	IMG_DATA[1303] = 32'h38708F;
	IMG_DATA[1304] = 32'h566065;
	IMG_DATA[1305] = 32'h969A91;
	IMG_DATA[1306] = 32'hC7C6B2;
	IMG_DATA[1307] = 32'hD1D0BD;
	IMG_DATA[1308] = 32'hABAA9A;
	IMG_DATA[1309] = 32'h3B4B5C;
	IMG_DATA[1310] = 32'h12375C;
	IMG_DATA[1311] = 32'h3A5972;
	IMG_DATA[1312] = 32'h64696D;
	IMG_DATA[1313] = 32'h5F6663;
	IMG_DATA[1314] = 32'h3B5B6F;
	IMG_DATA[1315] = 32'h50616D;
	IMG_DATA[1316] = 32'h92704C;
	IMG_DATA[1317] = 32'h926F4C;
	IMG_DATA[1318] = 32'h906D4B;
	IMG_DATA[1319] = 32'h906E4B;
	IMG_DATA[1320] = 32'h8F6F48;
	IMG_DATA[1321] = 32'h93704C;
	IMG_DATA[1322] = 32'h93704D;
	IMG_DATA[1323] = 32'h64584D;
	IMG_DATA[1324] = 32'h3A8BB2;
	IMG_DATA[1325] = 32'h5EC8EC;
	IMG_DATA[1326] = 32'h6FD2F5;
	IMG_DATA[1327] = 32'h77D5F6;
	IMG_DATA[1328] = 32'h80D6F6;
	IMG_DATA[1329] = 32'h92D9F8;
	IMG_DATA[1330] = 32'h9FDCF6;
	IMG_DATA[1331] = 32'h6CB0D2;
	IMG_DATA[1332] = 32'h5B83A4;
	IMG_DATA[1333] = 32'h62798F;
	IMG_DATA[1334] = 32'h6E7478;
	IMG_DATA[1335] = 32'h6D7371;
	IMG_DATA[1336] = 32'h3D5B6F;
	IMG_DATA[1337] = 32'h286083;
	IMG_DATA[1338] = 32'h30739B;
	IMG_DATA[1339] = 32'h447DA2;
	IMG_DATA[1340] = 32'h886949;
	IMG_DATA[1341] = 32'h8A6746;
	IMG_DATA[1342] = 32'h896846;
	IMG_DATA[1343] = 32'h896745;
	IMG_DATA[1344] = 32'h9F7B53;
	IMG_DATA[1345] = 32'h997851;
	IMG_DATA[1346] = 32'h94A1A5;
	IMG_DATA[1347] = 32'h81D3F4;
	IMG_DATA[1348] = 32'h84D9F8;
	IMG_DATA[1349] = 32'h88DAF9;
	IMG_DATA[1350] = 32'h8CD8F9;
	IMG_DATA[1351] = 32'h91D9F8;
	IMG_DATA[1352] = 32'h93D9F7;
	IMG_DATA[1353] = 32'h91D8F6;
	IMG_DATA[1354] = 32'h7ED1F3;
	IMG_DATA[1355] = 32'h6ECBEF;
	IMG_DATA[1356] = 32'h66C4E7;
	IMG_DATA[1357] = 32'h5CBADF;
	IMG_DATA[1358] = 32'h51AED3;
	IMG_DATA[1359] = 32'h4298BD;
	IMG_DATA[1360] = 32'h637377;
	IMG_DATA[1361] = 32'h9E7D53;
	IMG_DATA[1362] = 32'hA17F56;
	IMG_DATA[1363] = 32'h9C7D55;
	IMG_DATA[1364] = 32'h987C59;
	IMG_DATA[1365] = 32'h64ABC5;
	IMG_DATA[1366] = 32'h55B0D2;
	IMG_DATA[1367] = 32'h42A3CC;
	IMG_DATA[1368] = 32'h3386B4;
	IMG_DATA[1369] = 32'h355D7A;
	IMG_DATA[1370] = 32'h384C5F;
	IMG_DATA[1371] = 32'h384959;
	IMG_DATA[1372] = 32'h183E5D;
	IMG_DATA[1373] = 32'h27668D;
	IMG_DATA[1374] = 32'h42A0C9;
	IMG_DATA[1375] = 32'h43A6CF;
	IMG_DATA[1376] = 32'h357EAA;
	IMG_DATA[1377] = 32'h28658A;
	IMG_DATA[1378] = 32'h2D6086;
	IMG_DATA[1379] = 32'h426177;
	IMG_DATA[1380] = 32'h92714E;
	IMG_DATA[1381] = 32'h95734F;
	IMG_DATA[1382] = 32'h957450;
	IMG_DATA[1383] = 32'h94754E;
	IMG_DATA[1384] = 32'h95724D;
	IMG_DATA[1385] = 32'h93714C;
	IMG_DATA[1386] = 32'h886E55;
	IMG_DATA[1387] = 32'h4B515E;
	IMG_DATA[1388] = 32'h3E92BC;
	IMG_DATA[1389] = 32'h5BC6EB;
	IMG_DATA[1390] = 32'h6CD1F5;
	IMG_DATA[1391] = 32'h78D4F6;
	IMG_DATA[1392] = 32'h85D7F8;
	IMG_DATA[1393] = 32'h8AD7F7;
	IMG_DATA[1394] = 32'h94D8F7;
	IMG_DATA[1395] = 32'h8BD4F2;
	IMG_DATA[1396] = 32'h5CB3D7;
	IMG_DATA[1397] = 32'h317BA3;
	IMG_DATA[1398] = 32'h225A80;
	IMG_DATA[1399] = 32'h215B80;
	IMG_DATA[1400] = 32'h27698C;
	IMG_DATA[1401] = 32'h307AA1;
	IMG_DATA[1402] = 32'h3A8CB5;
	IMG_DATA[1403] = 32'h438CB8;
	IMG_DATA[1404] = 32'h866E55;
	IMG_DATA[1405] = 32'h8C6948;
	IMG_DATA[1406] = 32'h8B6948;
	IMG_DATA[1407] = 32'h8A6847;
	IMG_DATA[1408] = 32'hA28359;
	IMG_DATA[1409] = 32'hA28158;
	IMG_DATA[1410] = 32'h979893;
	IMG_DATA[1411] = 32'h80D0F4;
	IMG_DATA[1412] = 32'h84D7F7;
	IMG_DATA[1413] = 32'h87DAF8;
	IMG_DATA[1414] = 32'h8AD8F7;
	IMG_DATA[1415] = 32'h8CD9F8;
	IMG_DATA[1416] = 32'h91D9F9;
	IMG_DATA[1417] = 32'h92DAF5;
	IMG_DATA[1418] = 32'h84D5F4;
	IMG_DATA[1419] = 32'h71CEF0;
	IMG_DATA[1420] = 32'h66C6E9;
	IMG_DATA[1421] = 32'h5DBADF;
	IMG_DATA[1422] = 32'h51AFD4;
	IMG_DATA[1423] = 32'h439BBF;
	IMG_DATA[1424] = 32'h587583;
	IMG_DATA[1425] = 32'h9C7D54;
	IMG_DATA[1426] = 32'hA38058;
	IMG_DATA[1427] = 32'h9F7D53;
	IMG_DATA[1428] = 32'h9E7E58;
	IMG_DATA[1429] = 32'h5F9DB1;
	IMG_DATA[1430] = 32'h4CA7CC;
	IMG_DATA[1431] = 32'h46A9D3;
	IMG_DATA[1432] = 32'h42ACD8;
	IMG_DATA[1433] = 32'h3EA3D0;
	IMG_DATA[1434] = 32'h3C92BC;
	IMG_DATA[1435] = 32'h3F91B6;
	IMG_DATA[1436] = 32'h51A1C4;
	IMG_DATA[1437] = 32'h69BEDF;
	IMG_DATA[1438] = 32'h67C5E9;
	IMG_DATA[1439] = 32'h61C2E6;
	IMG_DATA[1440] = 32'h54B6DD;
	IMG_DATA[1441] = 32'h439DC4;
	IMG_DATA[1442] = 32'h3C85AA;
	IMG_DATA[1443] = 32'h3A6887;
	IMG_DATA[1444] = 32'h8A6F51;
	IMG_DATA[1445] = 32'h997851;
	IMG_DATA[1446] = 32'h977650;
	IMG_DATA[1447] = 32'h94744E;
	IMG_DATA[1448] = 32'h95734E;
	IMG_DATA[1449] = 32'h95724E;
	IMG_DATA[1450] = 32'h6B6158;
	IMG_DATA[1451] = 32'h354053;
	IMG_DATA[1452] = 32'h34799D;
	IMG_DATA[1453] = 32'h55C2E9;
	IMG_DATA[1454] = 32'h67CFF3;
	IMG_DATA[1455] = 32'h79D5F6;
	IMG_DATA[1456] = 32'h86D6F7;
	IMG_DATA[1457] = 32'h8CD6F6;
	IMG_DATA[1458] = 32'h8DD6F7;
	IMG_DATA[1459] = 32'h83D2F2;
	IMG_DATA[1460] = 32'h70C9EC;
	IMG_DATA[1461] = 32'h5DB7DD;
	IMG_DATA[1462] = 32'h4AA8CF;
	IMG_DATA[1463] = 32'h429DC3;
	IMG_DATA[1464] = 32'h419CC2;
	IMG_DATA[1465] = 32'h429EC6;
	IMG_DATA[1466] = 32'h44A0C8;
	IMG_DATA[1467] = 32'h4599C5;
	IMG_DATA[1468] = 32'h7F7467;
	IMG_DATA[1469] = 32'h92704E;
	IMG_DATA[1470] = 32'h8F6E4A;
	IMG_DATA[1471] = 32'h8D6C49;
	IMG_DATA[1472] = 32'hA5855C;
	IMG_DATA[1473] = 32'hA8875C;
	IMG_DATA[1474] = 32'h9E9688;
	IMG_DATA[1475] = 32'h7ED0F2;
	IMG_DATA[1476] = 32'h83D6F7;
	IMG_DATA[1477] = 32'h88D9F8;
	IMG_DATA[1478] = 32'h8BD8F8;
	IMG_DATA[1479] = 32'h8CD8F8;
	IMG_DATA[1480] = 32'h8DD8F8;
	IMG_DATA[1481] = 32'h91D9F7;
	IMG_DATA[1482] = 32'h87D6F4;
	IMG_DATA[1483] = 32'h70CEF0;
	IMG_DATA[1484] = 32'h63C5E8;
	IMG_DATA[1485] = 32'h5AB8DD;
	IMG_DATA[1486] = 32'h53AFD3;
	IMG_DATA[1487] = 32'h46A0C3;
	IMG_DATA[1488] = 32'h4F7B8F;
	IMG_DATA[1489] = 32'hA38258;
	IMG_DATA[1490] = 32'h9F7E55;
	IMG_DATA[1491] = 32'hA08056;
	IMG_DATA[1492] = 32'h997B53;
	IMG_DATA[1493] = 32'h465550;
	IMG_DATA[1494] = 32'h489FC3;
	IMG_DATA[1495] = 32'h46ABD3;
	IMG_DATA[1496] = 32'h44B3DC;
	IMG_DATA[1497] = 32'h4AB7DE;
	IMG_DATA[1498] = 32'h55B9E0;
	IMG_DATA[1499] = 32'h62BEE2;
	IMG_DATA[1500] = 32'h6AC5E7;
	IMG_DATA[1501] = 32'h73C7EA;
	IMG_DATA[1502] = 32'h68C2E7;
	IMG_DATA[1503] = 32'h64C1E6;
	IMG_DATA[1504] = 32'h60C0E6;
	IMG_DATA[1505] = 32'h54B5DB;
	IMG_DATA[1506] = 32'h469EC3;
	IMG_DATA[1507] = 32'h3C6F8C;
	IMG_DATA[1508] = 32'h725D40;
	IMG_DATA[1509] = 32'h987650;
	IMG_DATA[1510] = 32'h97754F;
	IMG_DATA[1511] = 32'h977450;
	IMG_DATA[1512] = 32'h987650;
	IMG_DATA[1513] = 32'h967350;
	IMG_DATA[1514] = 32'h4F4F56;
	IMG_DATA[1515] = 32'h293347;
	IMG_DATA[1516] = 32'h2D6284;
	IMG_DATA[1517] = 32'h4FBDE6;
	IMG_DATA[1518] = 32'h65CEF2;
	IMG_DATA[1519] = 32'h76D4F6;
	IMG_DATA[1520] = 32'h86D7F7;
	IMG_DATA[1521] = 32'h89D7F7;
	IMG_DATA[1522] = 32'h8CD6F7;
	IMG_DATA[1523] = 32'h81D2F5;
	IMG_DATA[1524] = 32'h7AD0F1;
	IMG_DATA[1525] = 32'h77CDEF;
	IMG_DATA[1526] = 32'h63C5E8;
	IMG_DATA[1527] = 32'h56BADF;
	IMG_DATA[1528] = 32'h53B2DA;
	IMG_DATA[1529] = 32'h50B1D9;
	IMG_DATA[1530] = 32'h4DABD7;
	IMG_DATA[1531] = 32'h4DA3D0;
	IMG_DATA[1532] = 32'h757978;
	IMG_DATA[1533] = 32'h93714D;
	IMG_DATA[1534] = 32'h95734E;
	IMG_DATA[1535] = 32'h906E4B;
	IMG_DATA[1536] = 32'hA5845B;
	IMG_DATA[1537] = 32'hA3835A;
	IMG_DATA[1538] = 32'h9C8A77;
	IMG_DATA[1539] = 32'h7CCDEF;
	IMG_DATA[1540] = 32'h80D6F7;
	IMG_DATA[1541] = 32'h89D9F9;
	IMG_DATA[1542] = 32'h8CDAFA;
	IMG_DATA[1543] = 32'h89D9F9;
	IMG_DATA[1544] = 32'h88D8F8;
	IMG_DATA[1545] = 32'h94D9F9;
	IMG_DATA[1546] = 32'h91DAF8;
	IMG_DATA[1547] = 32'h72CDF0;
	IMG_DATA[1548] = 32'h63C1E4;
	IMG_DATA[1549] = 32'h59B6DA;
	IMG_DATA[1550] = 32'h55B1D6;
	IMG_DATA[1551] = 32'h46A3C6;
	IMG_DATA[1552] = 32'h3F7A9A;
	IMG_DATA[1553] = 32'h605344;
	IMG_DATA[1554] = 32'h373531;
	IMG_DATA[1555] = 32'h363333;
	IMG_DATA[1556] = 32'h50453C;
	IMG_DATA[1557] = 32'h474534;
	IMG_DATA[1558] = 32'h4B5A57;
	IMG_DATA[1559] = 32'h45A4CD;
	IMG_DATA[1560] = 32'h46B5DE;
	IMG_DATA[1561] = 32'h50BCE3;
	IMG_DATA[1562] = 32'h61C3E9;
	IMG_DATA[1563] = 32'h6DCAED;
	IMG_DATA[1564] = 32'h5FAACC;
	IMG_DATA[1565] = 32'h152639;
	IMG_DATA[1566] = 32'h91323;
	IMG_DATA[1567] = 32'h5596B9;
	IMG_DATA[1568] = 32'h63C6EB;
	IMG_DATA[1569] = 32'h5CBDE5;
	IMG_DATA[1570] = 32'h4DA9D0;
	IMG_DATA[1571] = 32'h4A6065;
	IMG_DATA[1572] = 32'h635948;
	IMG_DATA[1573] = 32'h987650;
	IMG_DATA[1574] = 32'h997650;
	IMG_DATA[1575] = 32'h977650;
	IMG_DATA[1576] = 32'h997B53;
	IMG_DATA[1577] = 32'h8D7255;
	IMG_DATA[1578] = 32'h363F50;
	IMG_DATA[1579] = 32'h333E51;
	IMG_DATA[1580] = 32'h234D6C;
	IMG_DATA[1581] = 32'h4CB8E0;
	IMG_DATA[1582] = 32'h62CCEF;
	IMG_DATA[1583] = 32'h75D3F6;
	IMG_DATA[1584] = 32'h83D5F6;
	IMG_DATA[1585] = 32'h8DD6F7;
	IMG_DATA[1586] = 32'h87D5F5;
	IMG_DATA[1587] = 32'h7ED1F3;
	IMG_DATA[1588] = 32'h77CFF1;
	IMG_DATA[1589] = 32'h73CFF0;
	IMG_DATA[1590] = 32'h6DCAEC;
	IMG_DATA[1591] = 32'h66C3E7;
	IMG_DATA[1592] = 32'h5EBFE3;
	IMG_DATA[1593] = 32'h5BBCE3;
	IMG_DATA[1594] = 32'h56B7E0;
	IMG_DATA[1595] = 32'h4FA9D6;
	IMG_DATA[1596] = 32'h54768A;
	IMG_DATA[1597] = 32'h896D51;
	IMG_DATA[1598] = 32'h94724F;
	IMG_DATA[1599] = 32'h93714E;
	IMG_DATA[1600] = 32'hA5845C;
	IMG_DATA[1601] = 32'hA3835B;
	IMG_DATA[1602] = 32'h9E866E;
	IMG_DATA[1603] = 32'h7CCCEF;
	IMG_DATA[1604] = 32'h81D6F8;
	IMG_DATA[1605] = 32'h8BD9FA;
	IMG_DATA[1606] = 32'h8CDAFA;
	IMG_DATA[1607] = 32'h8BD9F8;
	IMG_DATA[1608] = 32'h87D6F6;
	IMG_DATA[1609] = 32'h8AD8F8;
	IMG_DATA[1610] = 32'h8AD9F7;
	IMG_DATA[1611] = 32'h6ECBED;
	IMG_DATA[1612] = 32'h5CB6DB;
	IMG_DATA[1613] = 32'h5CB5DB;
	IMG_DATA[1614] = 32'h5BB7DB;
	IMG_DATA[1615] = 32'h4AA7CB;
	IMG_DATA[1616] = 32'h367EA0;
	IMG_DATA[1617] = 32'h13212C;
	IMG_DATA[1618] = 32'h101922;
	IMG_DATA[1619] = 32'h101A27;
	IMG_DATA[1620] = 32'h18273F;
	IMG_DATA[1621] = 32'h1E3652;
	IMG_DATA[1622] = 32'h464A3E;
	IMG_DATA[1623] = 32'h525C56;
	IMG_DATA[1624] = 32'h45AAD3;
	IMG_DATA[1625] = 32'h54C1E7;
	IMG_DATA[1626] = 32'h67C8EB;
	IMG_DATA[1627] = 32'h81D1F2;
	IMG_DATA[1628] = 32'h8BCAE7;
	IMG_DATA[1629] = 32'h72A2BE;
	IMG_DATA[1630] = 32'h70B4D4;
	IMG_DATA[1631] = 32'h70C8ED;
	IMG_DATA[1632] = 32'h66C8EB;
	IMG_DATA[1633] = 32'h5ABBDF;
	IMG_DATA[1634] = 32'h5899B2;
	IMG_DATA[1635] = 32'h524C3D;
	IMG_DATA[1636] = 32'h495A65;
	IMG_DATA[1637] = 32'h93744E;
	IMG_DATA[1638] = 32'h977550;
	IMG_DATA[1639] = 32'h9A7652;
	IMG_DATA[1640] = 32'h9C7853;
	IMG_DATA[1641] = 32'h7A6755;
	IMG_DATA[1642] = 32'h3D495D;
	IMG_DATA[1643] = 32'h424D61;
	IMG_DATA[1644] = 32'h374A55;
	IMG_DATA[1645] = 32'h53AFD0;
	IMG_DATA[1646] = 32'h60C9EF;
	IMG_DATA[1647] = 32'h72D1F4;
	IMG_DATA[1648] = 32'h81D5F6;
	IMG_DATA[1649] = 32'h8ED6F6;
	IMG_DATA[1650] = 32'h8DD6F7;
	IMG_DATA[1651] = 32'h72B3CD;
	IMG_DATA[1652] = 32'h638591;
	IMG_DATA[1653] = 32'h6D8F9A;
	IMG_DATA[1654] = 32'h3D5E74;
	IMG_DATA[1655] = 32'h3B5D72;
	IMG_DATA[1656] = 32'h29506C;
	IMG_DATA[1657] = 32'h62BEE4;
	IMG_DATA[1658] = 32'h5ABCE3;
	IMG_DATA[1659] = 32'h4BAAD8;
	IMG_DATA[1660] = 32'h48677A;
	IMG_DATA[1661] = 32'h444245;
	IMG_DATA[1662] = 32'h977351;
	IMG_DATA[1663] = 32'h95714F;
	IMG_DATA[1664] = 32'hA8875B;
	IMG_DATA[1665] = 32'hA7865E;
	IMG_DATA[1666] = 32'hA18565;
	IMG_DATA[1667] = 32'h7AC7EA;
	IMG_DATA[1668] = 32'h80D6F6;
	IMG_DATA[1669] = 32'h8ADAF9;
	IMG_DATA[1670] = 32'h8BDAF9;
	IMG_DATA[1671] = 32'h8FDAF9;
	IMG_DATA[1672] = 32'h9ADCFA;
	IMG_DATA[1673] = 32'h95DAF9;
	IMG_DATA[1674] = 32'h80CFF1;
	IMG_DATA[1675] = 32'h6AC6E9;
	IMG_DATA[1676] = 32'h61C0E5;
	IMG_DATA[1677] = 32'h61C0E3;
	IMG_DATA[1678] = 32'h5AB7DA;
	IMG_DATA[1679] = 32'h4CA9CD;
	IMG_DATA[1680] = 32'h3982A6;
	IMG_DATA[1681] = 32'h142530;
	IMG_DATA[1682] = 32'hD141E;
	IMG_DATA[1683] = 32'h132033;
	IMG_DATA[1684] = 32'h243754;
	IMG_DATA[1685] = 32'h233959;
	IMG_DATA[1686] = 32'h317197;
	IMG_DATA[1687] = 32'h51594C;
	IMG_DATA[1688] = 32'h656D63;
	IMG_DATA[1689] = 32'h55B0D2;
	IMG_DATA[1690] = 32'h6EC0DE;
	IMG_DATA[1691] = 32'h83C2D7;
	IMG_DATA[1692] = 32'h93C3D0;
	IMG_DATA[1693] = 32'h95BEC4;
	IMG_DATA[1694] = 32'h87A9A7;
	IMG_DATA[1695] = 32'h8FA59B;
	IMG_DATA[1696] = 32'h858F7F;
	IMG_DATA[1697] = 32'h757562;
	IMG_DATA[1698] = 32'h71674E;
	IMG_DATA[1699] = 32'h495C64;
	IMG_DATA[1700] = 32'h3F6076;
	IMG_DATA[1701] = 32'h8C6A48;
	IMG_DATA[1702] = 32'h906C48;
	IMG_DATA[1703] = 32'h906D4C;
	IMG_DATA[1704] = 32'h97754F;
	IMG_DATA[1705] = 32'h6A5A4E;
	IMG_DATA[1706] = 32'h29354C;
	IMG_DATA[1707] = 32'h334055;
	IMG_DATA[1708] = 32'h464B55;
	IMG_DATA[1709] = 32'h79694B;
	IMG_DATA[1710] = 32'h749C9C;
	IMG_DATA[1711] = 32'h6CCEF3;
	IMG_DATA[1712] = 32'h7CD5F5;
	IMG_DATA[1713] = 32'h88D5F6;
	IMG_DATA[1714] = 32'h8DD7F7;
	IMG_DATA[1715] = 32'h27415B;
	IMG_DATA[1716] = 32'h3030B;
	IMG_DATA[1717] = 32'h2010B;
	IMG_DATA[1718] = 32'h20212;
	IMG_DATA[1719] = 32'h20211;
	IMG_DATA[1720] = 32'h11192D;
	IMG_DATA[1721] = 32'h67BDE1;
	IMG_DATA[1722] = 32'h58B9E4;
	IMG_DATA[1723] = 32'h47A0CE;
	IMG_DATA[1724] = 32'h444844;
	IMG_DATA[1725] = 32'h1A1B15;
	IMG_DATA[1726] = 32'h4A3E2A;
	IMG_DATA[1727] = 32'h94724F;
	IMG_DATA[1728] = 32'hA7875D;
	IMG_DATA[1729] = 32'hA9895D;
	IMG_DATA[1730] = 32'hA58765;
	IMG_DATA[1731] = 32'h79C2E5;
	IMG_DATA[1732] = 32'h7FD5F6;
	IMG_DATA[1733] = 32'h89D9F8;
	IMG_DATA[1734] = 32'h8CDAFA;
	IMG_DATA[1735] = 32'h8AD9F9;
	IMG_DATA[1736] = 32'h8EDAFA;
	IMG_DATA[1737] = 32'h8BD8F7;
	IMG_DATA[1738] = 32'h7DD4F5;
	IMG_DATA[1739] = 32'h6ECCEE;
	IMG_DATA[1740] = 32'h67C3E5;
	IMG_DATA[1741] = 32'h60BDE1;
	IMG_DATA[1742] = 32'h5BB5DA;
	IMG_DATA[1743] = 32'h4DA9CE;
	IMG_DATA[1744] = 32'h3985A8;
	IMG_DATA[1745] = 32'h202E37;
	IMG_DATA[1746] = 32'hD151F;
	IMG_DATA[1747] = 32'h1F2D3F;
	IMG_DATA[1748] = 32'h1E314E;
	IMG_DATA[1749] = 32'h192F4B;
	IMG_DATA[1750] = 32'h256A96;
	IMG_DATA[1751] = 32'h3A93BB;
	IMG_DATA[1752] = 32'h5E6655;
	IMG_DATA[1753] = 32'h5E563F;
	IMG_DATA[1754] = 32'h8D7C5B;
	IMG_DATA[1755] = 32'h8E7C54;
	IMG_DATA[1756] = 32'h8D784C;
	IMG_DATA[1757] = 32'h8F784A;
	IMG_DATA[1758] = 32'h887041;
	IMG_DATA[1759] = 32'h8B6F41;
	IMG_DATA[1760] = 32'h816437;
	IMG_DATA[1761] = 32'h6C5531;
	IMG_DATA[1762] = 32'h3C3930;
	IMG_DATA[1763] = 32'h3E738F;
	IMG_DATA[1764] = 32'h3F6076;
	IMG_DATA[1765] = 32'h80613F;
	IMG_DATA[1766] = 32'h8A6745;
	IMG_DATA[1767] = 32'h916D49;
	IMG_DATA[1768] = 32'h987450;
	IMG_DATA[1769] = 32'h6D5C4C;
	IMG_DATA[1770] = 32'h30394B;
	IMG_DATA[1771] = 32'h333D4F;
	IMG_DATA[1772] = 32'h2B3958;
	IMG_DATA[1773] = 32'h3F5B75;
	IMG_DATA[1774] = 32'h756E52;
	IMG_DATA[1775] = 32'h849F92;
	IMG_DATA[1776] = 32'h6FCEF1;
	IMG_DATA[1777] = 32'h7FD3F5;
	IMG_DATA[1778] = 32'h87D5F7;
	IMG_DATA[1779] = 32'h67ACCF;
	IMG_DATA[1780] = 32'h172941;
	IMG_DATA[1781] = 32'h10515;
	IMG_DATA[1782] = 32'hA132A;
	IMG_DATA[1783] = 32'h213957;
	IMG_DATA[1784] = 32'h65ABCE;
	IMG_DATA[1785] = 32'h62C1E9;
	IMG_DATA[1786] = 32'h56AAD4;
	IMG_DATA[1787] = 32'h5B8AA1;
	IMG_DATA[1788] = 32'h3D3428;
	IMG_DATA[1789] = 32'h1E211A;
	IMG_DATA[1790] = 32'h26261D;
	IMG_DATA[1791] = 32'h745A3D;
	IMG_DATA[1792] = 32'hA98A5E;
	IMG_DATA[1793] = 32'hA98A5F;
	IMG_DATA[1794] = 32'hA1865C;
	IMG_DATA[1795] = 32'h6DB9DC;
	IMG_DATA[1796] = 32'h81D5F8;
	IMG_DATA[1797] = 32'h8AD9F8;
	IMG_DATA[1798] = 32'h8BD9F9;
	IMG_DATA[1799] = 32'h8BD9F8;
	IMG_DATA[1800] = 32'h8AD8F9;
	IMG_DATA[1801] = 32'h84D7F7;
	IMG_DATA[1802] = 32'h7BD1F4;
	IMG_DATA[1803] = 32'h6ECBEE;
	IMG_DATA[1804] = 32'h66C4E5;
	IMG_DATA[1805] = 32'h62BDE1;
	IMG_DATA[1806] = 32'h5DB8DB;
	IMG_DATA[1807] = 32'h4EA9CC;
	IMG_DATA[1808] = 32'h4186A2;
	IMG_DATA[1809] = 32'h3E4140;
	IMG_DATA[1810] = 32'h11161C;
	IMG_DATA[1811] = 32'h252D32;
	IMG_DATA[1812] = 32'h1D2B42;
	IMG_DATA[1813] = 32'h1F385B;
	IMG_DATA[1814] = 32'h255E8B;
	IMG_DATA[1815] = 32'h3193C1;
	IMG_DATA[1816] = 32'h3F97BB;
	IMG_DATA[1817] = 32'h544835;
	IMG_DATA[1818] = 32'h7E6B48;
	IMG_DATA[1819] = 32'h8E7849;
	IMG_DATA[1820] = 32'h8D784C;
	IMG_DATA[1821] = 32'h887346;
	IMG_DATA[1822] = 32'h846C41;
	IMG_DATA[1823] = 32'h7D653C;
	IMG_DATA[1824] = 32'h7F6339;
	IMG_DATA[1825] = 32'h694E27;
	IMG_DATA[1826] = 32'h575547;
	IMG_DATA[1827] = 32'h417FA0;
	IMG_DATA[1828] = 32'h395B72;
	IMG_DATA[1829] = 32'h73553B;
	IMG_DATA[1830] = 32'h836340;
	IMG_DATA[1831] = 32'h8F6B49;
	IMG_DATA[1832] = 32'h987450;
	IMG_DATA[1833] = 32'h7B6349;
	IMG_DATA[1834] = 32'h242A37;
	IMG_DATA[1835] = 32'h2E3446;
	IMG_DATA[1836] = 32'h2E5168;
	IMG_DATA[1837] = 32'h2A3442;
	IMG_DATA[1838] = 32'h212624;
	IMG_DATA[1839] = 32'h7B6E4A;
	IMG_DATA[1840] = 32'h889B8C;
	IMG_DATA[1841] = 32'h74C7E6;
	IMG_DATA[1842] = 32'h7EC8E4;
	IMG_DATA[1843] = 32'h88CAE2;
	IMG_DATA[1844] = 32'h8BC6DB;
	IMG_DATA[1845] = 32'h88B6C7;
	IMG_DATA[1846] = 32'h88B3BD;
	IMG_DATA[1847] = 32'h82A4A6;
	IMG_DATA[1848] = 32'h83918B;
	IMG_DATA[1849] = 32'h787868;
	IMG_DATA[1850] = 32'h695E46;
	IMG_DATA[1851] = 32'h6A5A42;
	IMG_DATA[1852] = 32'h37302A;
	IMG_DATA[1853] = 32'h1B1914;
	IMG_DATA[1854] = 32'h221E14;
	IMG_DATA[1855] = 32'h614D33;
	IMG_DATA[1856] = 32'hAA8B60;
	IMG_DATA[1857] = 32'hAA895F;
	IMG_DATA[1858] = 32'h988051;
	IMG_DATA[1859] = 32'h6F9190;
	IMG_DATA[1860] = 32'h7BD4F5;
	IMG_DATA[1861] = 32'h86D9F8;
	IMG_DATA[1862] = 32'h89D9FA;
	IMG_DATA[1863] = 32'h8AD7F7;
	IMG_DATA[1864] = 32'h8AD6F7;
	IMG_DATA[1865] = 32'h83D6F5;
	IMG_DATA[1866] = 32'h7AD2F1;
	IMG_DATA[1867] = 32'h6ECBED;
	IMG_DATA[1868] = 32'h69C4E7;
	IMG_DATA[1869] = 32'h62BDE1;
	IMG_DATA[1870] = 32'h5DB7DA;
	IMG_DATA[1871] = 32'h4BA7C9;
	IMG_DATA[1872] = 32'h557B83;
	IMG_DATA[1873] = 32'h364C57;
	IMG_DATA[1874] = 32'h27343A;
	IMG_DATA[1875] = 32'hF0F0D;
	IMG_DATA[1876] = 32'h1B222D;
	IMG_DATA[1877] = 32'h30486D;
	IMG_DATA[1878] = 32'h1F456F;
	IMG_DATA[1879] = 32'h2982B2;
	IMG_DATA[1880] = 32'h3E9DC3;
	IMG_DATA[1881] = 32'h736140;
	IMG_DATA[1882] = 32'h82693E;
	IMG_DATA[1883] = 32'h8D7647;
	IMG_DATA[1884] = 32'h897348;
	IMG_DATA[1885] = 32'h937B4C;
	IMG_DATA[1886] = 32'h997F51;
	IMG_DATA[1887] = 32'h83673B;
	IMG_DATA[1888] = 32'h795B33;
	IMG_DATA[1889] = 32'h6D5029;
	IMG_DATA[1890] = 32'h615A48;
	IMG_DATA[1891] = 32'h3E7493;
	IMG_DATA[1892] = 32'h364A53;
	IMG_DATA[1893] = 32'h634A33;
	IMG_DATA[1894] = 32'h7B5C3C;
	IMG_DATA[1895] = 32'h876543;
	IMG_DATA[1896] = 32'h936F4C;
	IMG_DATA[1897] = 32'h947550;
	IMG_DATA[1898] = 32'h2C2D31;
	IMG_DATA[1899] = 32'h2A374A;
	IMG_DATA[1900] = 32'h3B6175;
	IMG_DATA[1901] = 32'h292A22;
	IMG_DATA[1902] = 32'h191A18;
	IMG_DATA[1903] = 32'h344A59;
	IMG_DATA[1904] = 32'h827856;
	IMG_DATA[1905] = 32'h736547;
	IMG_DATA[1906] = 32'h928766;
	IMG_DATA[1907] = 32'h958159;
	IMG_DATA[1908] = 32'h866F49;
	IMG_DATA[1909] = 32'h7E663D;
	IMG_DATA[1910] = 32'h7D663D;
	IMG_DATA[1911] = 32'h705630;
	IMG_DATA[1912] = 32'h725731;
	IMG_DATA[1913] = 32'h664D29;
	IMG_DATA[1914] = 32'h5E4827;
	IMG_DATA[1915] = 32'h44392D;
	IMG_DATA[1916] = 32'h4F4C4F;
	IMG_DATA[1917] = 32'h473D35;
	IMG_DATA[1918] = 32'h1B1710;
	IMG_DATA[1919] = 32'h362C1B;
	IMG_DATA[1920] = 32'hAD8E60;
	IMG_DATA[1921] = 32'hA8885F;
	IMG_DATA[1922] = 32'h98A7A7;
	IMG_DATA[1923] = 32'h82825F;
	IMG_DATA[1924] = 32'h75AFC5;
	IMG_DATA[1925] = 32'h84D7F7;
	IMG_DATA[1926] = 32'h8AD8F9;
	IMG_DATA[1927] = 32'h8AD8F8;
	IMG_DATA[1928] = 32'h85D6F6;
	IMG_DATA[1929] = 32'h7FD5F4;
	IMG_DATA[1930] = 32'h76D0F2;
	IMG_DATA[1931] = 32'h6FCBEC;
	IMG_DATA[1932] = 32'h64C4E5;
	IMG_DATA[1933] = 32'h63BCE0;
	IMG_DATA[1934] = 32'h5CB4D8;
	IMG_DATA[1935] = 32'h51A1C1;
	IMG_DATA[1936] = 32'h5F5F51;
	IMG_DATA[1937] = 32'h2E5066;
	IMG_DATA[1938] = 32'h386376;
	IMG_DATA[1939] = 32'h9090A;
	IMG_DATA[1940] = 32'h50606;
	IMG_DATA[1941] = 32'h151615;
	IMG_DATA[1942] = 32'hF1B2C;
	IMG_DATA[1943] = 32'h256A9C;
	IMG_DATA[1944] = 32'h3D8FB7;
	IMG_DATA[1945] = 32'h75603D;
	IMG_DATA[1946] = 32'h7B6237;
	IMG_DATA[1947] = 32'h856B3E;
	IMG_DATA[1948] = 32'h8E7649;
	IMG_DATA[1949] = 32'h927746;
	IMG_DATA[1950] = 32'h927344;
	IMG_DATA[1951] = 32'h88693D;
	IMG_DATA[1952] = 32'h785831;
	IMG_DATA[1953] = 32'h75542D;
	IMG_DATA[1954] = 32'h63553D;
	IMG_DATA[1955] = 32'h5A5C55;
	IMG_DATA[1956] = 32'h3C3B35;
	IMG_DATA[1957] = 32'h503C2B;
	IMG_DATA[1958] = 32'h77583B;
	IMG_DATA[1959] = 32'h916D48;
	IMG_DATA[1960] = 32'h9C7952;
	IMG_DATA[1961] = 32'h9F7C52;
	IMG_DATA[1962] = 32'h594734;
	IMG_DATA[1963] = 32'h2E5469;
	IMG_DATA[1964] = 32'h3D677B;
	IMG_DATA[1965] = 32'h222218;
	IMG_DATA[1966] = 32'h1F1D18;
	IMG_DATA[1967] = 32'h173F5B;
	IMG_DATA[1968] = 32'h549AB5;
	IMG_DATA[1969] = 32'h65563F;
	IMG_DATA[1970] = 32'h776644;
	IMG_DATA[1971] = 32'h8E7548;
	IMG_DATA[1972] = 32'h856C40;
	IMG_DATA[1973] = 32'h735C34;
	IMG_DATA[1974] = 32'h6C5630;
	IMG_DATA[1975] = 32'h66502D;
	IMG_DATA[1976] = 32'h664F2C;
	IMG_DATA[1977] = 32'h5F4826;
	IMG_DATA[1978] = 32'h594324;
	IMG_DATA[1979] = 32'h4C4332;
	IMG_DATA[1980] = 32'h535355;
	IMG_DATA[1981] = 32'h6E5946;
	IMG_DATA[1982] = 32'h1E2322;
	IMG_DATA[1983] = 32'h60533D;
	IMG_DATA[1984] = 32'hAB8D61;
	IMG_DATA[1985] = 32'hAA8C65;
	IMG_DATA[1986] = 32'h8BC2DA;
	IMG_DATA[1987] = 32'h6DB6C7;
	IMG_DATA[1988] = 32'h8A7D59;
	IMG_DATA[1989] = 32'h77B9CE;
	IMG_DATA[1990] = 32'h84D7F8;
	IMG_DATA[1991] = 32'h83D7F7;
	IMG_DATA[1992] = 32'h7ED5F5;
	IMG_DATA[1993] = 32'h7BD2F3;
	IMG_DATA[1994] = 32'h72CDEF;
	IMG_DATA[1995] = 32'h6BC8EB;
	IMG_DATA[1996] = 32'h64BFE1;
	IMG_DATA[1997] = 32'h63AFC9;
	IMG_DATA[1998] = 32'h5F909C;
	IMG_DATA[1999] = 32'h686D61;
	IMG_DATA[2000] = 32'h4E5148;
	IMG_DATA[2001] = 32'h193B60;
	IMG_DATA[2002] = 32'h3D7C9D;
	IMG_DATA[2003] = 32'h242625;
	IMG_DATA[2004] = 32'h221B14;
	IMG_DATA[2005] = 32'h110E0A;
	IMG_DATA[2006] = 32'h2F2416;
	IMG_DATA[2007] = 32'h3E413D;
	IMG_DATA[2008] = 32'h4C676F;
	IMG_DATA[2009] = 32'h796240;
	IMG_DATA[2010] = 32'h83653B;
	IMG_DATA[2011] = 32'h8D6E43;
	IMG_DATA[2012] = 32'h80673E;
	IMG_DATA[2013] = 32'h85673B;
	IMG_DATA[2014] = 32'h806137;
	IMG_DATA[2015] = 32'h7D5F39;
	IMG_DATA[2016] = 32'h7B5A30;
	IMG_DATA[2017] = 32'h75552D;
	IMG_DATA[2018] = 32'h654D2C;
	IMG_DATA[2019] = 32'h49341D;
	IMG_DATA[2020] = 32'h281F11;
	IMG_DATA[2021] = 32'h4A3625;
	IMG_DATA[2022] = 32'h7A5B3C;
	IMG_DATA[2023] = 32'h926E4B;
	IMG_DATA[2024] = 32'h9D7B52;
	IMG_DATA[2025] = 32'h997852;
	IMG_DATA[2026] = 32'h6A5340;
	IMG_DATA[2027] = 32'h40677F;
	IMG_DATA[2028] = 32'h242726;
	IMG_DATA[2029] = 32'h1F1B12;
	IMG_DATA[2030] = 32'hF1827;
	IMG_DATA[2031] = 32'h215C83;
	IMG_DATA[2032] = 32'h58AED3;
	IMG_DATA[2033] = 32'h847551;
	IMG_DATA[2034] = 32'h816B41;
	IMG_DATA[2035] = 32'h836C40;
	IMG_DATA[2036] = 32'h7E643A;
	IMG_DATA[2037] = 32'h816943;
	IMG_DATA[2038] = 32'h7E653E;
	IMG_DATA[2039] = 32'h785E38;
	IMG_DATA[2040] = 32'h674C2C;
	IMG_DATA[2041] = 32'h604828;
	IMG_DATA[2042] = 32'h533D20;
	IMG_DATA[2043] = 32'h514B38;
	IMG_DATA[2044] = 32'h625A51;
	IMG_DATA[2045] = 32'h886A4B;
	IMG_DATA[2046] = 32'h4E5759;
	IMG_DATA[2047] = 32'h807257;
	IMG_DATA[2048] = 32'hAB8D61;
	IMG_DATA[2049] = 32'hAA957A;
	IMG_DATA[2050] = 32'h86D1F3;
	IMG_DATA[2051] = 32'h4CB0E2;
	IMG_DATA[2052] = 32'h85B8BA;
	IMG_DATA[2053] = 32'h928059;
	IMG_DATA[2054] = 32'h829C96;
	IMG_DATA[2055] = 32'h8DAEAD;
	IMG_DATA[2056] = 32'h8BB4B7;
	IMG_DATA[2057] = 32'h88ACAE;
	IMG_DATA[2058] = 32'h8BA6A2;
	IMG_DATA[2059] = 32'h828F80;
	IMG_DATA[2060] = 32'h88826A;
	IMG_DATA[2061] = 32'h756245;
	IMG_DATA[2062] = 32'h654B2E;
	IMG_DATA[2063] = 32'h3B2C1D;
	IMG_DATA[2064] = 32'h3F6577;
	IMG_DATA[2065] = 32'h233F5C;
	IMG_DATA[2066] = 32'h316C95;
	IMG_DATA[2067] = 32'h435353;
	IMG_DATA[2068] = 32'h423221;
	IMG_DATA[2069] = 32'h433223;
	IMG_DATA[2070] = 32'h423020;
	IMG_DATA[2071] = 32'h3B2C1C;
	IMG_DATA[2072] = 32'h524029;
	IMG_DATA[2073] = 32'h6D5531;
	IMG_DATA[2074] = 32'h81633A;
	IMG_DATA[2075] = 32'h846438;
	IMG_DATA[2076] = 32'h78592F;
	IMG_DATA[2077] = 32'h76572E;
	IMG_DATA[2078] = 32'h6C4D28;
	IMG_DATA[2079] = 32'h6D4C26;
	IMG_DATA[2080] = 32'h75532E;
	IMG_DATA[2081] = 32'h694826;
	IMG_DATA[2082] = 32'h593F22;
	IMG_DATA[2083] = 32'h302416;
	IMG_DATA[2084] = 32'h201911;
	IMG_DATA[2085] = 32'h4E3827;
	IMG_DATA[2086] = 32'h846343;
	IMG_DATA[2087] = 32'h987551;
	IMG_DATA[2088] = 32'h9C7952;
	IMG_DATA[2089] = 32'h957F60;
	IMG_DATA[2090] = 32'h576371;
	IMG_DATA[2091] = 32'h54A3C9;
	IMG_DATA[2092] = 32'h23302F;
	IMG_DATA[2093] = 32'h161614;
	IMG_DATA[2094] = 32'h14324F;
	IMG_DATA[2095] = 32'h3581AC;
	IMG_DATA[2096] = 32'h5CACCE;
	IMG_DATA[2097] = 32'h87754F;
	IMG_DATA[2098] = 32'h7F653A;
	IMG_DATA[2099] = 32'h71582F;
	IMG_DATA[2100] = 32'h735932;
	IMG_DATA[2101] = 32'h795F39;
	IMG_DATA[2102] = 32'h7B5E35;
	IMG_DATA[2103] = 32'h7C5E39;
	IMG_DATA[2104] = 32'h664A2B;
	IMG_DATA[2105] = 32'h5E4527;
	IMG_DATA[2106] = 32'h573D22;
	IMG_DATA[2107] = 32'h514A3C;
	IMG_DATA[2108] = 32'h5A4F40;
	IMG_DATA[2109] = 32'h846546;
	IMG_DATA[2110] = 32'h92704D;
	IMG_DATA[2111] = 32'h997551;
	IMG_DATA[2112] = 32'hAD8F62;
	IMG_DATA[2113] = 32'hA59E92;
	IMG_DATA[2114] = 32'h7CD0F5;
	IMG_DATA[2115] = 32'h41A9E1;
	IMG_DATA[2116] = 32'h73D0F3;
	IMG_DATA[2117] = 32'h85ADA7;
	IMG_DATA[2118] = 32'h604B34;
	IMG_DATA[2119] = 32'h8B754B;
	IMG_DATA[2120] = 32'h8A7143;
	IMG_DATA[2121] = 32'h84683A;
	IMG_DATA[2122] = 32'h7D6033;
	IMG_DATA[2123] = 32'h795B30;
	IMG_DATA[2124] = 32'h77582F;
	IMG_DATA[2125] = 32'h6C4E28;
	IMG_DATA[2126] = 32'h654927;
	IMG_DATA[2127] = 32'h58422C;
	IMG_DATA[2128] = 32'h3D7590;
	IMG_DATA[2129] = 32'h2F4E62;
	IMG_DATA[2130] = 32'h265B85;
	IMG_DATA[2131] = 32'h456871;
	IMG_DATA[2132] = 32'h3E3021;
	IMG_DATA[2133] = 32'h3E2F21;
	IMG_DATA[2134] = 32'h3F2F21;
	IMG_DATA[2135] = 32'h3F3222;
	IMG_DATA[2136] = 32'h40301C;
	IMG_DATA[2137] = 32'h644A2A;
	IMG_DATA[2138] = 32'h624524;
	IMG_DATA[2139] = 32'h694926;
	IMG_DATA[2140] = 32'h684725;
	IMG_DATA[2141] = 32'h6C4D2C;
	IMG_DATA[2142] = 32'h6B4A28;
	IMG_DATA[2143] = 32'h5E3F21;
	IMG_DATA[2144] = 32'h573A1E;
	IMG_DATA[2145] = 32'h402A17;
	IMG_DATA[2146] = 32'h2B1D12;
	IMG_DATA[2147] = 32'h110D0B;
	IMG_DATA[2148] = 32'h261C16;
	IMG_DATA[2149] = 32'h60452F;
	IMG_DATA[2150] = 32'h8E6C48;
	IMG_DATA[2151] = 32'h9B7951;
	IMG_DATA[2152] = 32'h947651;
	IMG_DATA[2153] = 32'h41443F;
	IMG_DATA[2154] = 32'h2B383D;
	IMG_DATA[2155] = 32'h559EBF;
	IMG_DATA[2156] = 32'h395B68;
	IMG_DATA[2157] = 32'h1D1711;
	IMG_DATA[2158] = 32'h263B4B;
	IMG_DATA[2159] = 32'h418FB9;
	IMG_DATA[2160] = 32'h5DA5C3;
	IMG_DATA[2161] = 32'h806944;
	IMG_DATA[2162] = 32'h7B6037;
	IMG_DATA[2163] = 32'h765932;
	IMG_DATA[2164] = 32'h6E542F;
	IMG_DATA[2165] = 32'h755B38;
	IMG_DATA[2166] = 32'h6C502D;
	IMG_DATA[2167] = 32'h654A27;
	IMG_DATA[2168] = 32'h604829;
	IMG_DATA[2169] = 32'h5B4124;
	IMG_DATA[2170] = 32'h573E22;
	IMG_DATA[2171] = 32'h483B28;
	IMG_DATA[2172] = 32'h4D3E2A;
	IMG_DATA[2173] = 32'h785B3E;
	IMG_DATA[2174] = 32'h856746;
	IMG_DATA[2175] = 32'h8D6C4A;
	IMG_DATA[2176] = 32'hAC8C60;
	IMG_DATA[2177] = 32'h9EA19D;
	IMG_DATA[2178] = 32'h6FCCF2;
	IMG_DATA[2179] = 32'h429DD8;
	IMG_DATA[2180] = 32'h72CEF1;
	IMG_DATA[2181] = 32'h85D0E7;
	IMG_DATA[2182] = 32'h7F6B42;
	IMG_DATA[2183] = 32'h967B50;
	IMG_DATA[2184] = 32'h927745;
	IMG_DATA[2185] = 32'h7E6235;
	IMG_DATA[2186] = 32'h795D32;
	IMG_DATA[2187] = 32'h72562E;
	IMG_DATA[2188] = 32'h705730;
	IMG_DATA[2189] = 32'h664B29;
	IMG_DATA[2190] = 32'h5F4322;
	IMG_DATA[2191] = 32'h5D452C;
	IMG_DATA[2192] = 32'h41768F;
	IMG_DATA[2193] = 32'h274859;
	IMG_DATA[2194] = 32'h224567;
	IMG_DATA[2195] = 32'h41778B;
	IMG_DATA[2196] = 32'h3C2D20;
	IMG_DATA[2197] = 32'h3C2E21;
	IMG_DATA[2198] = 32'h3F2F20;
	IMG_DATA[2199] = 32'h423021;
	IMG_DATA[2200] = 32'h3B2B1D;
	IMG_DATA[2201] = 32'h332417;
	IMG_DATA[2202] = 32'h312011;
	IMG_DATA[2203] = 32'h332111;
	IMG_DATA[2204] = 32'h352212;
	IMG_DATA[2205] = 32'h332012;
	IMG_DATA[2206] = 32'h2D1E0F;
	IMG_DATA[2207] = 32'h23150C;
	IMG_DATA[2208] = 32'h1A110A;
	IMG_DATA[2209] = 32'h110B0A;
	IMG_DATA[2210] = 32'hC0707;
	IMG_DATA[2211] = 32'h18100E;
	IMG_DATA[2212] = 32'h4B3625;
	IMG_DATA[2213] = 32'h876442;
	IMG_DATA[2214] = 32'h97724C;
	IMG_DATA[2215] = 32'h94704A;
	IMG_DATA[2216] = 32'h7B5F41;
	IMG_DATA[2217] = 32'h39362B;
	IMG_DATA[2218] = 32'h2B2E2D;
	IMG_DATA[2219] = 32'h232727;
	IMG_DATA[2220] = 32'h1C1B18;
	IMG_DATA[2221] = 32'h312314;
	IMG_DATA[2222] = 32'h625136;
	IMG_DATA[2223] = 32'h7B7055;
	IMG_DATA[2224] = 32'h697568;
	IMG_DATA[2225] = 32'h836B43;
	IMG_DATA[2226] = 32'h785E35;
	IMG_DATA[2227] = 32'h775B34;
	IMG_DATA[2228] = 32'h6C512C;
	IMG_DATA[2229] = 32'h5F4729;
	IMG_DATA[2230] = 32'h5B4529;
	IMG_DATA[2231] = 32'h564026;
	IMG_DATA[2232] = 32'h543C23;
	IMG_DATA[2233] = 32'h593E22;
	IMG_DATA[2234] = 32'h563E23;
	IMG_DATA[2235] = 32'h42301A;
	IMG_DATA[2236] = 32'h453421;
	IMG_DATA[2237] = 32'h684D35;
	IMG_DATA[2238] = 32'h7B5C40;
	IMG_DATA[2239] = 32'h896745;
	IMG_DATA[2240] = 32'hAA8A5E;
	IMG_DATA[2241] = 32'h9CA2A2;
	IMG_DATA[2242] = 32'h6DC8F1;
	IMG_DATA[2243] = 32'h468DBF;
	IMG_DATA[2244] = 32'h6BCBF0;
	IMG_DATA[2245] = 32'h84D1EA;
	IMG_DATA[2246] = 32'h968251;
	IMG_DATA[2247] = 32'h957746;
	IMG_DATA[2248] = 32'h937544;
	IMG_DATA[2249] = 32'h90764C;
	IMG_DATA[2250] = 32'h846D41;
	IMG_DATA[2251] = 32'h81673F;
	IMG_DATA[2252] = 32'h715632;
	IMG_DATA[2253] = 32'h664D2A;
	IMG_DATA[2254] = 32'h5F4323;
	IMG_DATA[2255] = 32'h694F2F;
	IMG_DATA[2256] = 32'h3F6A7E;
	IMG_DATA[2257] = 32'h364345;
	IMG_DATA[2258] = 32'h23354B;
	IMG_DATA[2259] = 32'h4283A3;
	IMG_DATA[2260] = 32'h382C1F;
	IMG_DATA[2261] = 32'h493223;
	IMG_DATA[2262] = 32'h593E29;
	IMG_DATA[2263] = 32'h674B30;
	IMG_DATA[2264] = 32'h543A26;
	IMG_DATA[2265] = 32'h422D20;
	IMG_DATA[2266] = 32'h21170F;
	IMG_DATA[2267] = 32'h140F0B;
	IMG_DATA[2268] = 32'h90705;
	IMG_DATA[2269] = 32'hD0706;
	IMG_DATA[2270] = 32'hA0605;
	IMG_DATA[2271] = 32'hB0806;
	IMG_DATA[2272] = 32'h160E0A;
	IMG_DATA[2273] = 32'h291A12;
	IMG_DATA[2274] = 32'h432D1E;
	IMG_DATA[2275] = 32'h684A30;
	IMG_DATA[2276] = 32'h896642;
	IMG_DATA[2277] = 32'h946F4A;
	IMG_DATA[2278] = 32'h97724B;
	IMG_DATA[2279] = 32'h93704A;
	IMG_DATA[2280] = 32'h866644;
	IMG_DATA[2281] = 32'h4E3C27;
	IMG_DATA[2282] = 32'h4C412C;
	IMG_DATA[2283] = 32'h1B1714;
	IMG_DATA[2284] = 32'h191411;
	IMG_DATA[2285] = 32'h342515;
	IMG_DATA[2286] = 32'h6B5434;
	IMG_DATA[2287] = 32'h725833;
	IMG_DATA[2288] = 32'h75613F;
	IMG_DATA[2289] = 32'h705630;
	IMG_DATA[2290] = 32'h785C34;
	IMG_DATA[2291] = 32'h735731;
	IMG_DATA[2292] = 32'h664B29;
	IMG_DATA[2293] = 32'h5F4225;
	IMG_DATA[2294] = 32'h614727;
	IMG_DATA[2295] = 32'h553B21;
	IMG_DATA[2296] = 32'h553B20;
	IMG_DATA[2297] = 32'h553B20;
	IMG_DATA[2298] = 32'h543B21;
	IMG_DATA[2299] = 32'h3E2E1C;
	IMG_DATA[2300] = 32'h392D1E;
	IMG_DATA[2301] = 32'h634933;
	IMG_DATA[2302] = 32'h7F6042;
	IMG_DATA[2303] = 32'h8E6946;
	IMG_DATA[2304] = 32'hAB8B5F;
	IMG_DATA[2305] = 32'h98A2A3;
	IMG_DATA[2306] = 32'h68C2E6;
	IMG_DATA[2307] = 32'h446476;
	IMG_DATA[2308] = 32'h5DBEE6;
	IMG_DATA[2309] = 32'h7ECDE8;
	IMG_DATA[2310] = 32'h988254;
	IMG_DATA[2311] = 32'h8C6E3B;
	IMG_DATA[2312] = 32'h886C3D;
	IMG_DATA[2313] = 32'h8B7044;
	IMG_DATA[2314] = 32'h8F6F41;
	IMG_DATA[2315] = 32'h917042;
	IMG_DATA[2316] = 32'h72542D;
	IMG_DATA[2317] = 32'h664A2A;
	IMG_DATA[2318] = 32'h644824;
	IMG_DATA[2319] = 32'h5F4728;
	IMG_DATA[2320] = 32'h4C473B;
	IMG_DATA[2321] = 32'h473925;
	IMG_DATA[2322] = 32'h16181F;
	IMG_DATA[2323] = 32'h295577;
	IMG_DATA[2324] = 32'h2B251F;
	IMG_DATA[2325] = 32'h4E3724;
	IMG_DATA[2326] = 32'h68492E;
	IMG_DATA[2327] = 32'h805C3C;
	IMG_DATA[2328] = 32'h886440;
	IMG_DATA[2329] = 32'h856240;
	IMG_DATA[2330] = 32'h704F33;
	IMG_DATA[2331] = 32'h4C3422;
	IMG_DATA[2332] = 32'h422F1E;
	IMG_DATA[2333] = 32'h593E29;
	IMG_DATA[2334] = 32'h593E28;
	IMG_DATA[2335] = 32'h513925;
	IMG_DATA[2336] = 32'h6D4E32;
	IMG_DATA[2337] = 32'h835F3D;
	IMG_DATA[2338] = 32'h926C47;
	IMG_DATA[2339] = 32'h97734C;
	IMG_DATA[2340] = 32'h9A754F;
	IMG_DATA[2341] = 32'h97724C;
	IMG_DATA[2342] = 32'h946F49;
	IMG_DATA[2343] = 32'h98744D;
	IMG_DATA[2344] = 32'h95734C;
	IMG_DATA[2345] = 32'h715538;
	IMG_DATA[2346] = 32'h3A291B;
	IMG_DATA[2347] = 32'h1D1610;
	IMG_DATA[2348] = 32'h18120D;
	IMG_DATA[2349] = 32'h31241A;
	IMG_DATA[2350] = 32'h382C1C;
	IMG_DATA[2351] = 32'h59452C;
	IMG_DATA[2352] = 32'h6E5739;
	IMG_DATA[2353] = 32'h7B5E38;
	IMG_DATA[2354] = 32'h694D2B;
	IMG_DATA[2355] = 32'h614525;
	IMG_DATA[2356] = 32'h614426;
	IMG_DATA[2357] = 32'h5C3F23;
	IMG_DATA[2358] = 32'h634A2D;
	IMG_DATA[2359] = 32'h563B22;
	IMG_DATA[2360] = 32'h52381E;
	IMG_DATA[2361] = 32'h4A331D;
	IMG_DATA[2362] = 32'h382714;
	IMG_DATA[2363] = 32'h312518;
	IMG_DATA[2364] = 32'h403123;
	IMG_DATA[2365] = 32'h5B432D;
	IMG_DATA[2366] = 32'h7E5E3F;
	IMG_DATA[2367] = 32'h8B6643;
	IMG_DATA[2368] = 32'hA8885C;
	IMG_DATA[2369] = 32'h97A3A3;
	IMG_DATA[2370] = 32'h61B8D9;
	IMG_DATA[2371] = 32'h625C44;
	IMG_DATA[2372] = 32'h8B9686;
	IMG_DATA[2373] = 32'h76AEBC;
	IMG_DATA[2374] = 32'h98855B;
	IMG_DATA[2375] = 32'h927642;
	IMG_DATA[2376] = 32'h8C6E3F;
	IMG_DATA[2377] = 32'h84693F;
	IMG_DATA[2378] = 32'h816134;
	IMG_DATA[2379] = 32'h7A5931;
	IMG_DATA[2380] = 32'h6D512D;
	IMG_DATA[2381] = 32'h644926;
	IMG_DATA[2382] = 32'h6B4D29;
	IMG_DATA[2383] = 32'h654A29;
	IMG_DATA[2384] = 32'h4A3822;
	IMG_DATA[2385] = 32'h3F2F1B;
	IMG_DATA[2386] = 32'h1D150F;
	IMG_DATA[2387] = 32'h14100A;
	IMG_DATA[2388] = 32'h251C12;
	IMG_DATA[2389] = 32'h4B3522;
	IMG_DATA[2390] = 32'h6F5032;
	IMG_DATA[2391] = 32'h85603E;
	IMG_DATA[2392] = 32'h9A754E;
	IMG_DATA[2393] = 32'h9A744E;
	IMG_DATA[2394] = 32'h96714A;
	IMG_DATA[2395] = 32'h97724C;
	IMG_DATA[2396] = 32'h936D47;
	IMG_DATA[2397] = 32'h936E48;
	IMG_DATA[2398] = 32'h916C47;
	IMG_DATA[2399] = 32'h936E48;
	IMG_DATA[2400] = 32'h97714B;
	IMG_DATA[2401] = 32'h96714B;
	IMG_DATA[2402] = 32'h9A744E;
	IMG_DATA[2403] = 32'h9B764F;
	IMG_DATA[2404] = 32'h99764F;
	IMG_DATA[2405] = 32'h96714B;
	IMG_DATA[2406] = 32'h946F49;
	IMG_DATA[2407] = 32'h97714C;
	IMG_DATA[2408] = 32'h96714B;
	IMG_DATA[2409] = 32'h9C7750;
	IMG_DATA[2410] = 32'h98734C;
	IMG_DATA[2411] = 32'h765637;
	IMG_DATA[2412] = 32'h5B422B;
	IMG_DATA[2413] = 32'h443020;
	IMG_DATA[2414] = 32'h322518;
	IMG_DATA[2415] = 32'h281C12;
	IMG_DATA[2416] = 32'h362514;
	IMG_DATA[2417] = 32'h452F1A;
	IMG_DATA[2418] = 32'h49331C;
	IMG_DATA[2419] = 32'h49331B;
	IMG_DATA[2420] = 32'h452F19;
	IMG_DATA[2421] = 32'h412D19;
	IMG_DATA[2422] = 32'h412F1B;
	IMG_DATA[2423] = 32'h392815;
	IMG_DATA[2424] = 32'h302112;
	IMG_DATA[2425] = 32'h271C11;
	IMG_DATA[2426] = 32'h221914;
	IMG_DATA[2427] = 32'h2E241A;
	IMG_DATA[2428] = 32'h5B422C;
	IMG_DATA[2429] = 32'h755639;
	IMG_DATA[2430] = 32'h7E5D3C;
	IMG_DATA[2431] = 32'h896441;
	IMG_DATA[2432] = 32'hAA8C5F;
	IMG_DATA[2433] = 32'h899DA4;
	IMG_DATA[2434] = 32'h59AACD;
	IMG_DATA[2435] = 32'h6D593F;
	IMG_DATA[2436] = 32'h998256;
	IMG_DATA[2437] = 32'h977E51;
	IMG_DATA[2438] = 32'h91784B;
	IMG_DATA[2439] = 32'h907343;
	IMG_DATA[2440] = 32'h8B6D3D;
	IMG_DATA[2441] = 32'h7A5C34;
	IMG_DATA[2442] = 32'h6C502C;
	IMG_DATA[2443] = 32'h634729;
	IMG_DATA[2444] = 32'h5D4223;
	IMG_DATA[2445] = 32'h624623;
	IMG_DATA[2446] = 32'h644827;
	IMG_DATA[2447] = 32'h5E4122;
	IMG_DATA[2448] = 32'h493520;
	IMG_DATA[2449] = 32'h291E11;
	IMG_DATA[2450] = 32'h90504;
	IMG_DATA[2451] = 32'h140E09;
	IMG_DATA[2452] = 32'h1E170F;
	IMG_DATA[2453] = 32'h493322;
	IMG_DATA[2454] = 32'h755639;
	IMG_DATA[2455] = 32'h936F49;
	IMG_DATA[2456] = 32'h99744D;
	IMG_DATA[2457] = 32'h99734E;
	IMG_DATA[2458] = 32'h9B7650;
	IMG_DATA[2459] = 32'h9A754F;
	IMG_DATA[2460] = 32'h98734D;
	IMG_DATA[2461] = 32'h96714B;
	IMG_DATA[2462] = 32'h96714B;
	IMG_DATA[2463] = 32'h9A7650;
	IMG_DATA[2464] = 32'h98734C;
	IMG_DATA[2465] = 32'h9C7850;
	IMG_DATA[2466] = 32'h9C7750;
	IMG_DATA[2467] = 32'h9E7A53;
	IMG_DATA[2468] = 32'h9D7850;
	IMG_DATA[2469] = 32'h9B7750;
	IMG_DATA[2470] = 32'h97724C;
	IMG_DATA[2471] = 32'h9A754F;
	IMG_DATA[2472] = 32'h9C784F;
	IMG_DATA[2473] = 32'h9C7850;
	IMG_DATA[2474] = 32'h9A7650;
	IMG_DATA[2475] = 32'h8A6643;
	IMG_DATA[2476] = 32'h745437;
	IMG_DATA[2477] = 32'h63472E;
	IMG_DATA[2478] = 32'h473222;
	IMG_DATA[2479] = 32'h33251A;
	IMG_DATA[2480] = 32'h1C140F;
	IMG_DATA[2481] = 32'h1D140C;
	IMG_DATA[2482] = 32'h1B120A;
	IMG_DATA[2483] = 32'h180E08;
	IMG_DATA[2484] = 32'h130C07;
	IMG_DATA[2485] = 32'h130C06;
	IMG_DATA[2486] = 32'h130D07;
	IMG_DATA[2487] = 32'h1A120E;
	IMG_DATA[2488] = 32'h1E1512;
	IMG_DATA[2489] = 32'h221815;
	IMG_DATA[2490] = 32'h281D17;
	IMG_DATA[2491] = 32'h4A3523;
	IMG_DATA[2492] = 32'h7E5B3B;
	IMG_DATA[2493] = 32'h8D6843;
	IMG_DATA[2494] = 32'h8C6641;
	IMG_DATA[2495] = 32'h906A46;
	IMG_DATA[2496] = 32'hA8895E;
	IMG_DATA[2497] = 32'h4E5149;
	IMG_DATA[2498] = 32'h324A52;
	IMG_DATA[2499] = 32'h5E4933;
	IMG_DATA[2500] = 32'h846A45;
	IMG_DATA[2501] = 32'h856C45;
	IMG_DATA[2502] = 32'h977A4C;
	IMG_DATA[2503] = 32'h87673A;
	IMG_DATA[2504] = 32'h7D5D32;
	IMG_DATA[2505] = 32'h72532B;
	IMG_DATA[2506] = 32'h6C4D28;
	IMG_DATA[2507] = 32'h6B4E2C;
	IMG_DATA[2508] = 32'h5D4121;
	IMG_DATA[2509] = 32'h5D4222;
	IMG_DATA[2510] = 32'h51381E;
	IMG_DATA[2511] = 32'h3E2815;
	IMG_DATA[2512] = 32'h312113;
	IMG_DATA[2513] = 32'h221812;
	IMG_DATA[2514] = 32'hB0805;
	IMG_DATA[2515] = 32'h150F09;
	IMG_DATA[2516] = 32'h261D15;
	IMG_DATA[2517] = 32'h3B2B1E;
	IMG_DATA[2518] = 32'h7F5F3F;
	IMG_DATA[2519] = 32'h99754E;
	IMG_DATA[2520] = 32'h9A754F;
	IMG_DATA[2521] = 32'h97724C;
	IMG_DATA[2522] = 32'h99744F;
	IMG_DATA[2523] = 32'h98734E;
	IMG_DATA[2524] = 32'h946F49;
	IMG_DATA[2525] = 32'h97724C;
	IMG_DATA[2526] = 32'h97724C;
	IMG_DATA[2527] = 32'h9A754F;
	IMG_DATA[2528] = 32'h9B7750;
	IMG_DATA[2529] = 32'h9D7851;
	IMG_DATA[2530] = 32'h9E7A51;
	IMG_DATA[2531] = 32'h9E7B51;
	IMG_DATA[2532] = 32'h9B7750;
	IMG_DATA[2533] = 32'h9A754E;
	IMG_DATA[2534] = 32'h9A754F;
	IMG_DATA[2535] = 32'h9C7650;
	IMG_DATA[2536] = 32'h9B774E;
	IMG_DATA[2537] = 32'h99744D;
	IMG_DATA[2538] = 32'h9A744F;
	IMG_DATA[2539] = 32'h95704A;
	IMG_DATA[2540] = 32'h8D6A45;
	IMG_DATA[2541] = 32'h866341;
	IMG_DATA[2542] = 32'h705134;
	IMG_DATA[2543] = 32'h553C28;
	IMG_DATA[2544] = 32'h3E2D1E;
	IMG_DATA[2545] = 32'h130C0A;
	IMG_DATA[2546] = 32'h40201;
	IMG_DATA[2547] = 32'h110C07;
	IMG_DATA[2548] = 32'h140E0A;
	IMG_DATA[2549] = 32'h80504;
	IMG_DATA[2550] = 32'h30201;
	IMG_DATA[2551] = 32'h80706;
	IMG_DATA[2552] = 32'h2E2119;
	IMG_DATA[2553] = 32'h483222;
	IMG_DATA[2554] = 32'h61442E;
	IMG_DATA[2555] = 32'h7F5C3C;
	IMG_DATA[2556] = 32'h8C6542;
	IMG_DATA[2557] = 32'h88643F;
	IMG_DATA[2558] = 32'h8E6A42;
	IMG_DATA[2559] = 32'h906944;
	IMG_DATA[2560] = 32'hA28158;
	IMG_DATA[2561] = 32'h4D442A;
	IMG_DATA[2562] = 32'h252318;
	IMG_DATA[2563] = 32'h56402E;
	IMG_DATA[2564] = 32'h94754C;
	IMG_DATA[2565] = 32'h684D2D;
	IMG_DATA[2566] = 32'h755532;
	IMG_DATA[2567] = 32'h684A28;
	IMG_DATA[2568] = 32'h604323;
	IMG_DATA[2569] = 32'h5A3E21;
	IMG_DATA[2570] = 32'h54391D;
	IMG_DATA[2571] = 32'h533A22;
	IMG_DATA[2572] = 32'h442C16;
	IMG_DATA[2573] = 32'h392313;
	IMG_DATA[2574] = 32'h2F1F11;
	IMG_DATA[2575] = 32'h221811;
	IMG_DATA[2576] = 32'h1B1411;
	IMG_DATA[2577] = 32'h1D1413;
	IMG_DATA[2578] = 32'h17100F;
	IMG_DATA[2579] = 32'h1F1711;
	IMG_DATA[2580] = 32'h34281C;
	IMG_DATA[2581] = 32'h674D35;
	IMG_DATA[2582] = 32'h8F6B48;
	IMG_DATA[2583] = 32'h97724C;
	IMG_DATA[2584] = 32'h95724C;
	IMG_DATA[2585] = 32'h916C48;
	IMG_DATA[2586] = 32'h916E49;
	IMG_DATA[2587] = 32'h95704B;
	IMG_DATA[2588] = 32'h97734D;
	IMG_DATA[2589] = 32'h95724B;
	IMG_DATA[2590] = 32'h99744E;
	IMG_DATA[2591] = 32'h99744E;
	IMG_DATA[2592] = 32'h9A754E;
	IMG_DATA[2593] = 32'h9A764F;
	IMG_DATA[2594] = 32'h9C7750;
	IMG_DATA[2595] = 32'h9A764F;
	IMG_DATA[2596] = 32'h98754E;
	IMG_DATA[2597] = 32'h97724D;
	IMG_DATA[2598] = 32'h936F49;
	IMG_DATA[2599] = 32'h95704A;
	IMG_DATA[2600] = 32'h99744E;
	IMG_DATA[2601] = 32'h96714B;
	IMG_DATA[2602] = 32'h946E4A;
	IMG_DATA[2603] = 32'h946F49;
	IMG_DATA[2604] = 32'h906B46;
	IMG_DATA[2605] = 32'h906B45;
	IMG_DATA[2606] = 32'h8D6744;
	IMG_DATA[2607] = 32'h886441;
	IMG_DATA[2608] = 32'h6C4E33;
	IMG_DATA[2609] = 32'h1F1915;
	IMG_DATA[2610] = 32'h181410;
	IMG_DATA[2611] = 32'h3F2C1C;
	IMG_DATA[2612] = 32'h5D4029;
	IMG_DATA[2613] = 32'h513924;
	IMG_DATA[2614] = 32'h24190E;
	IMG_DATA[2615] = 32'h19150F;
	IMG_DATA[2616] = 32'h3C2B1B;
	IMG_DATA[2617] = 32'h835D3B;
	IMG_DATA[2618] = 32'h8B6440;
	IMG_DATA[2619] = 32'h916743;
	IMG_DATA[2620] = 32'h916843;
	IMG_DATA[2621] = 32'h8F6743;
	IMG_DATA[2622] = 32'h946C44;
	IMG_DATA[2623] = 32'h966E45;
	IMG_DATA[2624] = 32'hA28259;
	IMG_DATA[2625] = 32'h373120;
	IMG_DATA[2626] = 32'h29271C;
	IMG_DATA[2627] = 32'h1A170E;
	IMG_DATA[2628] = 32'h2D1E15;
	IMG_DATA[2629] = 32'h4C3724;
	IMG_DATA[2630] = 32'h402D1E;
	IMG_DATA[2631] = 32'h3C2919;
	IMG_DATA[2632] = 32'h332212;
	IMG_DATA[2633] = 32'h2D1D11;
	IMG_DATA[2634] = 32'h28190E;
	IMG_DATA[2635] = 32'h1C130C;
	IMG_DATA[2636] = 32'h1A0E09;
	IMG_DATA[2637] = 32'h1B1109;
	IMG_DATA[2638] = 32'h1D140E;
	IMG_DATA[2639] = 32'h140F0F;
	IMG_DATA[2640] = 32'h151010;
	IMG_DATA[2641] = 32'h1C1412;
	IMG_DATA[2642] = 32'h2B1F17;
	IMG_DATA[2643] = 32'h5E442D;
	IMG_DATA[2644] = 32'h806040;
	IMG_DATA[2645] = 32'h8F6D49;
	IMG_DATA[2646] = 32'h8D6A47;
	IMG_DATA[2647] = 32'h8E6C48;
	IMG_DATA[2648] = 32'h916D4A;
	IMG_DATA[2649] = 32'h93714B;
	IMG_DATA[2650] = 32'h93724C;
	IMG_DATA[2651] = 32'h95724D;
	IMG_DATA[2652] = 32'h96714C;
	IMG_DATA[2653] = 32'h94704A;
	IMG_DATA[2654] = 32'h96704B;
	IMG_DATA[2655] = 32'h96714C;
	IMG_DATA[2656] = 32'h97724C;
	IMG_DATA[2657] = 32'h95714B;
	IMG_DATA[2658] = 32'h96714B;
	IMG_DATA[2659] = 32'h95724B;
	IMG_DATA[2660] = 32'h95734B;
	IMG_DATA[2661] = 32'h9A754F;
	IMG_DATA[2662] = 32'h97724C;
	IMG_DATA[2663] = 32'h95704A;
	IMG_DATA[2664] = 32'h956F4A;
	IMG_DATA[2665] = 32'h96704A;
	IMG_DATA[2666] = 32'h906B45;
	IMG_DATA[2667] = 32'h8E6A45;
	IMG_DATA[2668] = 32'h8A6641;
	IMG_DATA[2669] = 32'h8B6541;
	IMG_DATA[2670] = 32'h8A6340;
	IMG_DATA[2671] = 32'h8D6543;
	IMG_DATA[2672] = 32'h845E3C;
	IMG_DATA[2673] = 32'h563E28;
	IMG_DATA[2674] = 32'h583E27;
	IMG_DATA[2675] = 32'h825D3C;
	IMG_DATA[2676] = 32'h8E6642;
	IMG_DATA[2677] = 32'h8D6440;
	IMG_DATA[2678] = 32'h89613D;
	IMG_DATA[2679] = 32'h7A5837;
	IMG_DATA[2680] = 32'h7F5B36;
	IMG_DATA[2681] = 32'h8E6740;
	IMG_DATA[2682] = 32'h8F6841;
	IMG_DATA[2683] = 32'h926842;
	IMG_DATA[2684] = 32'h956A44;
	IMG_DATA[2685] = 32'h987048;
	IMG_DATA[2686] = 32'h987045;
	IMG_DATA[2687] = 32'h9A7246;
	IMG_DATA[2688] = 32'h9D7951;
	IMG_DATA[2689] = 32'h4C3D24;
	IMG_DATA[2690] = 32'h252015;
	IMG_DATA[2691] = 32'h15110B;
	IMG_DATA[2692] = 32'h281F15;
	IMG_DATA[2693] = 32'h402F1F;
	IMG_DATA[2694] = 32'h563D28;
	IMG_DATA[2695] = 32'h4D3725;
	IMG_DATA[2696] = 32'h342619;
	IMG_DATA[2697] = 32'h16120D;
	IMG_DATA[2698] = 32'hB0806;
	IMG_DATA[2699] = 32'hB0706;
	IMG_DATA[2700] = 32'h60302;
	IMG_DATA[2701] = 32'h40202;
	IMG_DATA[2702] = 32'hA0708;
	IMG_DATA[2703] = 32'h1F1712;
	IMG_DATA[2704] = 32'h3C2C1D;
	IMG_DATA[2705] = 32'h59412C;
	IMG_DATA[2706] = 32'h715336;
	IMG_DATA[2707] = 32'h8A6743;
	IMG_DATA[2708] = 32'h916C49;
	IMG_DATA[2709] = 32'h8E6C49;
	IMG_DATA[2710] = 32'h936F4A;
	IMG_DATA[2711] = 32'h8E6A47;
	IMG_DATA[2712] = 32'h936F4A;
	IMG_DATA[2713] = 32'h94704A;
	IMG_DATA[2714] = 32'h8F6D48;
	IMG_DATA[2715] = 32'h93704C;
	IMG_DATA[2716] = 32'h95714C;
	IMG_DATA[2717] = 32'h8D6946;
	IMG_DATA[2718] = 32'h926E4A;
	IMG_DATA[2719] = 32'h916D48;
	IMG_DATA[2720] = 32'h926E48;
	IMG_DATA[2721] = 32'h946F49;
	IMG_DATA[2722] = 32'h916C46;
	IMG_DATA[2723] = 32'h95704A;
	IMG_DATA[2724] = 32'h96714B;
	IMG_DATA[2725] = 32'h95704A;
	IMG_DATA[2726] = 32'h926D47;
	IMG_DATA[2727] = 32'h8E6945;
	IMG_DATA[2728] = 32'h8C6842;
	IMG_DATA[2729] = 32'h8E6943;
	IMG_DATA[2730] = 32'h8C6742;
	IMG_DATA[2731] = 32'h8A6441;
	IMG_DATA[2732] = 32'h8F6944;
	IMG_DATA[2733] = 32'h936C44;
	IMG_DATA[2734] = 32'h8F6742;
	IMG_DATA[2735] = 32'h8C6440;
	IMG_DATA[2736] = 32'h89633D;
	IMG_DATA[2737] = 32'h8C643F;
	IMG_DATA[2738] = 32'h8E663E;
	IMG_DATA[2739] = 32'h946942;
	IMG_DATA[2740] = 32'h936943;
	IMG_DATA[2741] = 32'h946741;
	IMG_DATA[2742] = 32'h906641;
	IMG_DATA[2743] = 32'h906640;
	IMG_DATA[2744] = 32'h936A42;
	IMG_DATA[2745] = 32'h986D44;
	IMG_DATA[2746] = 32'h956D44;
	IMG_DATA[2747] = 32'h9B6F46;
	IMG_DATA[2748] = 32'h9C7047;
	IMG_DATA[2749] = 32'h9C7348;
	IMG_DATA[2750] = 32'h9F784C;
	IMG_DATA[2751] = 32'hA47A4E;
	IMG_DATA[2752] = 32'h99744D;
	IMG_DATA[2753] = 32'h9A7750;
	IMG_DATA[2754] = 32'h554229;
	IMG_DATA[2755] = 32'h261E14;
	IMG_DATA[2756] = 32'h3A2B1D;
	IMG_DATA[2757] = 32'h61472D;
	IMG_DATA[2758] = 32'h886642;
	IMG_DATA[2759] = 32'h725336;
	IMG_DATA[2760] = 32'h372B1E;
	IMG_DATA[2761] = 32'h90605;
	IMG_DATA[2762] = 32'hC0705;
	IMG_DATA[2763] = 32'h38261B;
	IMG_DATA[2764] = 32'h322317;
	IMG_DATA[2765] = 32'h16110C;
	IMG_DATA[2766] = 32'h1C1917;
	IMG_DATA[2767] = 32'h241C16;
	IMG_DATA[2768] = 32'h7D5C3D;
	IMG_DATA[2769] = 32'h936F49;
	IMG_DATA[2770] = 32'h926D48;
	IMG_DATA[2771] = 32'h946D49;
	IMG_DATA[2772] = 32'h906E4A;
	IMG_DATA[2773] = 32'h936E4A;
	IMG_DATA[2774] = 32'h916E4A;
	IMG_DATA[2775] = 32'h916E49;
	IMG_DATA[2776] = 32'h906D48;
	IMG_DATA[2777] = 32'h8E6A47;
	IMG_DATA[2778] = 32'h8C6A47;
	IMG_DATA[2779] = 32'h946E4A;
	IMG_DATA[2780] = 32'h906C48;
	IMG_DATA[2781] = 32'h866542;
	IMG_DATA[2782] = 32'h856442;
	IMG_DATA[2783] = 32'h886644;
	IMG_DATA[2784] = 32'h8A6643;
	IMG_DATA[2785] = 32'h926D49;
	IMG_DATA[2786] = 32'h906B45;
	IMG_DATA[2787] = 32'h906B45;
	IMG_DATA[2788] = 32'h916D46;
	IMG_DATA[2789] = 32'h906B46;
	IMG_DATA[2790] = 32'h906C46;
	IMG_DATA[2791] = 32'h886241;
	IMG_DATA[2792] = 32'h86613F;
	IMG_DATA[2793] = 32'h896341;
	IMG_DATA[2794] = 32'h86633F;
	IMG_DATA[2795] = 32'h86623F;
	IMG_DATA[2796] = 32'h8A6441;
	IMG_DATA[2797] = 32'h8D6741;
	IMG_DATA[2798] = 32'h8B6640;
	IMG_DATA[2799] = 32'h8E6841;
	IMG_DATA[2800] = 32'h926A44;
	IMG_DATA[2801] = 32'h986D44;
	IMG_DATA[2802] = 32'h976C44;
	IMG_DATA[2803] = 32'h926A41;
	IMG_DATA[2804] = 32'h91673F;
	IMG_DATA[2805] = 32'h926841;
	IMG_DATA[2806] = 32'h906740;
	IMG_DATA[2807] = 32'h8D653E;
	IMG_DATA[2808] = 32'h926841;
	IMG_DATA[2809] = 32'h926941;
	IMG_DATA[2810] = 32'h966D46;
	IMG_DATA[2811] = 32'h9A6F45;
	IMG_DATA[2812] = 32'h9F7348;
	IMG_DATA[2813] = 32'h9B7146;
	IMG_DATA[2814] = 32'h9F7549;
	IMG_DATA[2815] = 32'h9E7548;
	IMG_DATA[2816] = 32'h936F49;
	IMG_DATA[2817] = 32'h97734D;
	IMG_DATA[2818] = 32'h926F4A;
	IMG_DATA[2819] = 32'h715638;
	IMG_DATA[2820] = 32'h846242;
	IMG_DATA[2821] = 32'h946F49;
	IMG_DATA[2822] = 32'h926C46;
	IMG_DATA[2823] = 32'h8E6945;
	IMG_DATA[2824] = 32'h403526;
	IMG_DATA[2825] = 32'h201E19;
	IMG_DATA[2826] = 32'h332217;
	IMG_DATA[2827] = 32'h815D40;
	IMG_DATA[2828] = 32'h876340;
	IMG_DATA[2829] = 32'h6B5034;
	IMG_DATA[2830] = 32'h513D29;
	IMG_DATA[2831] = 32'h58402A;
	IMG_DATA[2832] = 32'h8F6B46;
	IMG_DATA[2833] = 32'h956F4B;
	IMG_DATA[2834] = 32'h926D49;
	IMG_DATA[2835] = 32'h96714C;
	IMG_DATA[2836] = 32'h926E48;
	IMG_DATA[2837] = 32'h906B46;
	IMG_DATA[2838] = 32'h916D49;
	IMG_DATA[2839] = 32'h8E6B48;
	IMG_DATA[2840] = 32'h8C6745;
	IMG_DATA[2841] = 32'h8E6945;
	IMG_DATA[2842] = 32'h8D6A48;
	IMG_DATA[2843] = 32'h8E6943;
	IMG_DATA[2844] = 32'h8F6A46;
	IMG_DATA[2845] = 32'h896945;
	IMG_DATA[2846] = 32'h856440;
	IMG_DATA[2847] = 32'h8A6643;
	IMG_DATA[2848] = 32'h8F6C46;
	IMG_DATA[2849] = 32'h8E6A43;
	IMG_DATA[2850] = 32'h8D6844;
	IMG_DATA[2851] = 32'h906C46;
	IMG_DATA[2852] = 32'h906B45;
	IMG_DATA[2853] = 32'h916D46;
	IMG_DATA[2854] = 32'h936C46;
	IMG_DATA[2855] = 32'h8D6842;
	IMG_DATA[2856] = 32'h8D6842;
	IMG_DATA[2857] = 32'h8A6541;
	IMG_DATA[2858] = 32'h84603D;
	IMG_DATA[2859] = 32'h825E3B;
	IMG_DATA[2860] = 32'h83603C;
	IMG_DATA[2861] = 32'h835E3A;
	IMG_DATA[2862] = 32'h8B653F;
	IMG_DATA[2863] = 32'h8F6841;
	IMG_DATA[2864] = 32'h976D45;
	IMG_DATA[2865] = 32'h9F764A;
	IMG_DATA[2866] = 32'h976D44;
	IMG_DATA[2867] = 32'h946942;
	IMG_DATA[2868] = 32'h92673F;
	IMG_DATA[2869] = 32'h906640;
	IMG_DATA[2870] = 32'h91683F;
	IMG_DATA[2871] = 32'h8F6740;
	IMG_DATA[2872] = 32'h916942;
	IMG_DATA[2873] = 32'h976D45;
	IMG_DATA[2874] = 32'h956A42;
	IMG_DATA[2875] = 32'h956A42;
	IMG_DATA[2876] = 32'h946B41;
	IMG_DATA[2877] = 32'h936C43;
	IMG_DATA[2878] = 32'h91683F;
	IMG_DATA[2879] = 32'h966D43;
	IMG_DATA[2880] = 32'h95714B;
	IMG_DATA[2881] = 32'h97724C;
	IMG_DATA[2882] = 32'h96714B;
	IMG_DATA[2883] = 32'h956F4A;
	IMG_DATA[2884] = 32'h97724C;
	IMG_DATA[2885] = 32'h96724B;
	IMG_DATA[2886] = 32'h95704A;
	IMG_DATA[2887] = 32'h95704A;
	IMG_DATA[2888] = 32'h725639;
	IMG_DATA[2889] = 32'h684E33;
	IMG_DATA[2890] = 32'h826041;
	IMG_DATA[2891] = 32'h926E48;
	IMG_DATA[2892] = 32'h936D49;
	IMG_DATA[2893] = 32'h946E4A;
	IMG_DATA[2894] = 32'h8F6B47;
	IMG_DATA[2895] = 32'h906B46;
	IMG_DATA[2896] = 32'h8C6741;
	IMG_DATA[2897] = 32'h8F6A46;
	IMG_DATA[2898] = 32'h926D48;
	IMG_DATA[2899] = 32'h8F6945;
	IMG_DATA[2900] = 32'h8E6945;
	IMG_DATA[2901] = 32'h8F6946;
	IMG_DATA[2902] = 32'h8C6843;
	IMG_DATA[2903] = 32'h8B6743;
	IMG_DATA[2904] = 32'h8D6845;
	IMG_DATA[2905] = 32'h8D6943;
	IMG_DATA[2906] = 32'h8D6943;
	IMG_DATA[2907] = 32'h8E6945;
	IMG_DATA[2908] = 32'h906B45;
	IMG_DATA[2909] = 32'h8A6741;
	IMG_DATA[2910] = 32'h8C6844;
	IMG_DATA[2911] = 32'h8B6744;
	IMG_DATA[2912] = 32'h886440;
	IMG_DATA[2913] = 32'h8A6641;
	IMG_DATA[2914] = 32'h8B6640;
	IMG_DATA[2915] = 32'h8D6643;
	IMG_DATA[2916] = 32'h8D6844;
	IMG_DATA[2917] = 32'h8B6640;
	IMG_DATA[2918] = 32'h906A43;
	IMG_DATA[2919] = 32'h916C44;
	IMG_DATA[2920] = 32'h8F6943;
	IMG_DATA[2921] = 32'h8A633F;
	IMG_DATA[2922] = 32'h89623F;
	IMG_DATA[2923] = 32'h815C3B;
	IMG_DATA[2924] = 32'h7F5A37;
	IMG_DATA[2925] = 32'h85603D;
	IMG_DATA[2926] = 32'h86613C;
	IMG_DATA[2927] = 32'h8B653E;
	IMG_DATA[2928] = 32'h926A42;
	IMG_DATA[2929] = 32'h946A42;
	IMG_DATA[2930] = 32'h90683F;
	IMG_DATA[2931] = 32'h91673F;
	IMG_DATA[2932] = 32'h9B7145;
	IMG_DATA[2933] = 32'h956D42;
	IMG_DATA[2934] = 32'h8C653E;
	IMG_DATA[2935] = 32'h8A633D;
	IMG_DATA[2936] = 32'h8B643D;
	IMG_DATA[2937] = 32'h845D38;
	IMG_DATA[2938] = 32'h8C633E;
	IMG_DATA[2939] = 32'h8D633D;
	IMG_DATA[2940] = 32'h8C633C;
	IMG_DATA[2941] = 32'h875E3A;
	IMG_DATA[2942] = 32'h8A613C;
	IMG_DATA[2943] = 32'h8F653D;
	IMG_DATA[2944] = 32'h8D6A47;
	IMG_DATA[2945] = 32'h906B48;
	IMG_DATA[2946] = 32'h916C47;
	IMG_DATA[2947] = 32'h936D49;
	IMG_DATA[2948] = 32'h96714B;
	IMG_DATA[2949] = 32'h95704A;
	IMG_DATA[2950] = 32'h98734D;
	IMG_DATA[2951] = 32'h98734D;
	IMG_DATA[2952] = 32'h9D784F;
	IMG_DATA[2953] = 32'h9C764F;
	IMG_DATA[2954] = 32'h99734E;
	IMG_DATA[2955] = 32'h96714B;
	IMG_DATA[2956] = 32'h926D47;
	IMG_DATA[2957] = 32'h8E6943;
	IMG_DATA[2958] = 32'h906B46;
	IMG_DATA[2959] = 32'h8E6943;
	IMG_DATA[2960] = 32'h8F6A45;
	IMG_DATA[2961] = 32'h8E6945;
	IMG_DATA[2962] = 32'h8E6946;
	IMG_DATA[2963] = 32'h8C6844;
	IMG_DATA[2964] = 32'h8E6845;
	IMG_DATA[2965] = 32'h8D6744;
	IMG_DATA[2966] = 32'h8B6740;
	IMG_DATA[2967] = 32'h8F6B45;
	IMG_DATA[2968] = 32'h8B6542;
	IMG_DATA[2969] = 32'h8F6A45;
	IMG_DATA[2970] = 32'h896542;
	IMG_DATA[2971] = 32'h896440;
	IMG_DATA[2972] = 32'h86603E;
	IMG_DATA[2973] = 32'h886440;
	IMG_DATA[2974] = 32'h8B6743;
	IMG_DATA[2975] = 32'h876440;
	IMG_DATA[2976] = 32'h88643D;
	IMG_DATA[2977] = 32'h896542;
	IMG_DATA[2978] = 32'h8B6542;
	IMG_DATA[2979] = 32'h8F6845;
	IMG_DATA[2980] = 32'h8B6540;
	IMG_DATA[2981] = 32'h896340;
	IMG_DATA[2982] = 32'h8A6540;
	IMG_DATA[2983] = 32'h8C6541;
	IMG_DATA[2984] = 32'h896340;
	IMG_DATA[2985] = 32'h89623F;
	IMG_DATA[2986] = 32'h8B6440;
	IMG_DATA[2987] = 32'h8D643F;
	IMG_DATA[2988] = 32'h855F3C;
	IMG_DATA[2989] = 32'h88613E;
	IMG_DATA[2990] = 32'h87613E;
	IMG_DATA[2991] = 32'h87623A;
	IMG_DATA[2992] = 32'h89623D;
	IMG_DATA[2993] = 32'h8F683E;
	IMG_DATA[2994] = 32'h8A613B;
	IMG_DATA[2995] = 32'h855E39;
	IMG_DATA[2996] = 32'h875E3A;
	IMG_DATA[2997] = 32'h8C633C;
	IMG_DATA[2998] = 32'h8E653C;
	IMG_DATA[2999] = 32'h855D35;
	IMG_DATA[3000] = 32'h815A35;
	IMG_DATA[3001] = 32'h7E5834;
	IMG_DATA[3002] = 32'h7F5734;
	IMG_DATA[3003] = 32'h7D5732;
	IMG_DATA[3004] = 32'h855B33;
	IMG_DATA[3005] = 32'h8A6039;
	IMG_DATA[3006] = 32'h845933;
	IMG_DATA[3007] = 32'h875D36;
	IMG_DATA[3008] = 32'h8A6845;
	IMG_DATA[3009] = 32'h8F6C4A;
	IMG_DATA[3010] = 32'h8E6B48;
	IMG_DATA[3011] = 32'h926D48;
	IMG_DATA[3012] = 32'h96714B;
	IMG_DATA[3013] = 32'h956F4A;
	IMG_DATA[3014] = 32'h99754D;
	IMG_DATA[3015] = 32'hA17951;
	IMG_DATA[3016] = 32'h9E7950;
	IMG_DATA[3017] = 32'hA07B52;
	IMG_DATA[3018] = 32'h9B764E;
	IMG_DATA[3019] = 32'h946F49;
	IMG_DATA[3020] = 32'h936E49;
	IMG_DATA[3021] = 32'h957049;
	IMG_DATA[3022] = 32'h8E6944;
	IMG_DATA[3023] = 32'h95704A;
	IMG_DATA[3024] = 32'h906A45;
	IMG_DATA[3025] = 32'h8D6743;
	IMG_DATA[3026] = 32'h8F6B46;
	IMG_DATA[3027] = 32'h926E48;
	IMG_DATA[3028] = 32'h8E6943;
	IMG_DATA[3029] = 32'h8B6643;
	IMG_DATA[3030] = 32'h8B6543;
	IMG_DATA[3031] = 32'h886441;
	IMG_DATA[3032] = 32'h896240;
	IMG_DATA[3033] = 32'h85603E;
	IMG_DATA[3034] = 32'h86623F;
	IMG_DATA[3035] = 32'h896541;
	IMG_DATA[3036] = 32'h87633D;
	IMG_DATA[3037] = 32'h896441;
	IMG_DATA[3038] = 32'h87623F;
	IMG_DATA[3039] = 32'h85603D;
	IMG_DATA[3040] = 32'h876240;
	IMG_DATA[3041] = 32'h8A6541;
	IMG_DATA[3042] = 32'h88633E;
	IMG_DATA[3043] = 32'h89633E;
	IMG_DATA[3044] = 32'h88633E;
	IMG_DATA[3045] = 32'h89613E;
	IMG_DATA[3046] = 32'h87603C;
	IMG_DATA[3047] = 32'h87613D;
	IMG_DATA[3048] = 32'h835E3C;
	IMG_DATA[3049] = 32'h7E5C39;
	IMG_DATA[3050] = 32'h845E3A;
	IMG_DATA[3051] = 32'h86603C;
	IMG_DATA[3052] = 32'h835C3B;
	IMG_DATA[3053] = 32'h7E5A37;
	IMG_DATA[3054] = 32'h7E5936;
	IMG_DATA[3055] = 32'h865F3A;
	IMG_DATA[3056] = 32'h805A38;
	IMG_DATA[3057] = 32'h7E5734;
	IMG_DATA[3058] = 32'h7A5634;
	IMG_DATA[3059] = 32'h775332;
	IMG_DATA[3060] = 32'h795332;
	IMG_DATA[3061] = 32'h734D2C;
	IMG_DATA[3062] = 32'h815933;
	IMG_DATA[3063] = 32'h875C34;
	IMG_DATA[3064] = 32'h845B33;
	IMG_DATA[3065] = 32'h835A33;
	IMG_DATA[3066] = 32'h896036;
	IMG_DATA[3067] = 32'h835933;
	IMG_DATA[3068] = 32'h7A512D;
	IMG_DATA[3069] = 32'h805832;
	IMG_DATA[3070] = 32'h815832;
	IMG_DATA[3071] = 32'h79512C;
end
